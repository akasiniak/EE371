module s2pShiftRegister;
endmodule
