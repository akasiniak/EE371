module johnsonCounter(count, clk, reset);
  input clk, reset;
  output [3:0] count;
endmodule
