module bitSampleCount;
endmodule
