module bitIdentifierCount;
endmodule
