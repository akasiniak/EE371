module startBitDetect;
endmodule
