module p2sShiftRegister;
endmodule
