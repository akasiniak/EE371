// Copyright (C) 2017  Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License 
// Subscription Agreement, the Intel Quartus Prime License Agreement,
// the Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is for
// the sole purpose of programming logic devices manufactured by
// Intel and sold by Intel or its authorized distributors.  Please
// refer to the applicable agreement for further details.

// VENDOR "Altera"
// PROGRAM "Quartus Prime"
// VERSION "Version 17.1.0 Build 590 10/25/2017 SJ Standard Edition"

// DATE "02/06/2018 13:42:06"

// 
// Device: Altera 5CSEMA5F31C6 Package FBGA896
// 

// 
// This greybox netlist file is for third party Synthesis Tools
// for timing and resource estimation only.
// 


module processor (
	altera_reserved_tms,
	altera_reserved_tck,
	altera_reserved_tdi,
	altera_reserved_tdo,
	clk_clk,
	led_pio_external_connection_export,
	reset_reset_n,
	switches_pio_external_connection_export)/* synthesis synthesis_greybox=1 */;
input 	altera_reserved_tms;
input 	altera_reserved_tck;
input 	altera_reserved_tdi;
output 	altera_reserved_tdo;
input 	clk_clk;
output 	[9:0] led_pio_external_connection_export;
input 	reset_reset_n;
input 	[9:0] switches_pio_external_connection_export;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \cpu|M_st_data[8]~q ;
wire \cpu|M_st_data[9]~q ;
wire \onchip_mem|the_altsyncram|auto_generated|q_a[0] ;
wire \onchip_mem|the_altsyncram|auto_generated|q_a[16] ;
wire \onchip_mem|the_altsyncram|auto_generated|q_a[8] ;
wire \onchip_mem|the_altsyncram|auto_generated|q_a[24] ;
wire \onchip_mem|the_altsyncram|auto_generated|q_a[5] ;
wire \onchip_mem|the_altsyncram|auto_generated|q_a[21] ;
wire \onchip_mem|the_altsyncram|auto_generated|q_a[13] ;
wire \onchip_mem|the_altsyncram|auto_generated|q_a[29] ;
wire \onchip_mem|the_altsyncram|auto_generated|q_a[4] ;
wire \onchip_mem|the_altsyncram|auto_generated|q_a[20] ;
wire \onchip_mem|the_altsyncram|auto_generated|q_a[12] ;
wire \onchip_mem|the_altsyncram|auto_generated|q_a[28] ;
wire \onchip_mem|the_altsyncram|auto_generated|q_a[6] ;
wire \onchip_mem|the_altsyncram|auto_generated|q_a[22] ;
wire \onchip_mem|the_altsyncram|auto_generated|q_a[14] ;
wire \onchip_mem|the_altsyncram|auto_generated|q_a[30] ;
wire \onchip_mem|the_altsyncram|auto_generated|q_a[7] ;
wire \onchip_mem|the_altsyncram|auto_generated|q_a[23] ;
wire \onchip_mem|the_altsyncram|auto_generated|q_a[15] ;
wire \onchip_mem|the_altsyncram|auto_generated|q_a[31] ;
wire \onchip_mem|the_altsyncram|auto_generated|q_a[11] ;
wire \onchip_mem|the_altsyncram|auto_generated|q_a[27] ;
wire \onchip_mem|the_altsyncram|auto_generated|q_a[10] ;
wire \onchip_mem|the_altsyncram|auto_generated|q_a[26] ;
wire \onchip_mem|the_altsyncram|auto_generated|q_a[25] ;
wire \onchip_mem|the_altsyncram|auto_generated|q_a[9] ;
wire \onchip_mem|the_altsyncram|auto_generated|q_a[3] ;
wire \onchip_mem|the_altsyncram|auto_generated|q_a[19] ;
wire \onchip_mem|the_altsyncram|auto_generated|q_a[2] ;
wire \onchip_mem|the_altsyncram|auto_generated|q_a[18] ;
wire \onchip_mem|the_altsyncram|auto_generated|q_a[1] ;
wire \onchip_mem|the_altsyncram|auto_generated|q_a[17] ;
wire \cpu|the_processor_cpu_nios2_oci|readdata[0]~q ;
wire \jtag_uart|the_processor_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[0] ;
wire \jtag_uart|Add1~1_sumout ;
wire \cpu|the_processor_cpu_nios2_oci|readdata[16]~q ;
wire \cpu|M_st_data[16]~q ;
wire \cpu|the_processor_cpu_nios2_oci|readdata[8]~q ;
wire \cpu|the_processor_cpu_nios2_oci|readdata[24]~q ;
wire \cpu|the_processor_cpu_nios2_oci|readdata[5]~q ;
wire \jtag_uart|the_processor_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[5] ;
wire \cpu|the_processor_cpu_nios2_oci|readdata[21]~q ;
wire \cpu|M_st_data[21]~q ;
wire \jtag_uart|Add1~5_sumout ;
wire \cpu|the_processor_cpu_nios2_oci|readdata[13]~q ;
wire \cpu|M_st_data[13]~q ;
wire \cpu|the_processor_cpu_nios2_oci|readdata[29]~q ;
wire \cpu|the_processor_cpu_nios2_oci|readdata[4]~q ;
wire \jtag_uart|the_processor_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[4] ;
wire \cpu|the_processor_cpu_nios2_oci|readdata[20]~q ;
wire \cpu|M_st_data[20]~q ;
wire \jtag_uart|Add1~9_sumout ;
wire \cpu|the_processor_cpu_nios2_oci|readdata[12]~q ;
wire \cpu|M_st_data[12]~q ;
wire \cpu|the_processor_cpu_nios2_oci|readdata[28]~q ;
wire \cpu|the_processor_cpu_nios2_oci|readdata[6]~q ;
wire \jtag_uart|the_processor_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[6] ;
wire \cpu|the_processor_cpu_nios2_oci|readdata[22]~q ;
wire \cpu|M_st_data[22]~q ;
wire \jtag_uart|Add1~13_sumout ;
wire \cpu|the_processor_cpu_nios2_oci|readdata[14]~q ;
wire \cpu|M_st_data[14]~q ;
wire \cpu|the_processor_cpu_nios2_oci|readdata[30]~q ;
wire \cpu|the_processor_cpu_nios2_oci|readdata[7]~q ;
wire \jtag_uart|the_processor_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[7] ;
wire \cpu|the_processor_cpu_nios2_oci|readdata[23]~q ;
wire \cpu|M_st_data[23]~q ;
wire \cpu|the_processor_cpu_nios2_oci|readdata[15]~q ;
wire \cpu|M_st_data[15]~q ;
wire \cpu|the_processor_cpu_nios2_oci|readdata[31]~q ;
wire \cpu|the_processor_cpu_nios2_oci|readdata[11]~q ;
wire \cpu|M_st_data[11]~q ;
wire \cpu|the_processor_cpu_nios2_oci|readdata[27]~q ;
wire \cpu|the_processor_cpu_nios2_oci|readdata[10]~q ;
wire \cpu|M_st_data[10]~q ;
wire \cpu|the_processor_cpu_nios2_oci|readdata[26]~q ;
wire \cpu|the_processor_cpu_nios2_oci|readdata[25]~q ;
wire \cpu|the_processor_cpu_nios2_oci|readdata[9]~q ;
wire \jtag_uart|the_processor_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[3] ;
wire \cpu|the_processor_cpu_nios2_oci|readdata[3]~q ;
wire \cpu|the_processor_cpu_nios2_oci|readdata[19]~q ;
wire \cpu|M_st_data[19]~q ;
wire \jtag_uart|Add1~17_sumout ;
wire \jtag_uart|the_processor_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[2] ;
wire \cpu|the_processor_cpu_nios2_oci|readdata[2]~q ;
wire \jtag_uart|Add1~21_sumout ;
wire \cpu|the_processor_cpu_nios2_oci|readdata[18]~q ;
wire \cpu|M_st_data[18]~q ;
wire \jtag_uart|the_processor_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[1] ;
wire \cpu|the_processor_cpu_nios2_oci|readdata[1]~q ;
wire \cpu|the_processor_cpu_nios2_oci|readdata[17]~q ;
wire \cpu|M_st_data[17]~q ;
wire \jtag_uart|Add1~25_sumout ;
wire \led_pio|data_out[0]~q ;
wire \led_pio|data_out[1]~q ;
wire \led_pio|data_out[2]~q ;
wire \led_pio|data_out[3]~q ;
wire \led_pio|data_out[4]~q ;
wire \led_pio|data_out[5]~q ;
wire \led_pio|data_out[6]~q ;
wire \led_pio|data_out[7]~q ;
wire \led_pio|data_out[8]~q ;
wire \led_pio|data_out[9]~q ;
wire \cpu|the_processor_cpu_nios2_oci|the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_tck|sr[0]~q ;
wire \cpu|the_processor_cpu_nios2_oci|the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_tck|ir_out[0]~q ;
wire \cpu|the_processor_cpu_nios2_oci|the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_tck|ir_out[1]~q ;
wire \jtag_uart|processor_jtag_uart_alt_jtag_atlantic|tdo~q ;
wire \cpu|M_st_data[0]~q ;
wire \rst_controller|r_sync_rst~q ;
wire \cpu|clr_break_line~q ;
wire \cpu|d_write~q ;
wire \mm_interconnect_0|led_pio_s1_agent_rsp_fifo|mem_used[1]~q ;
wire \cpu|M_alu_result[5]~q ;
wire \cpu|M_alu_result[4]~q ;
wire \cpu|M_alu_result[6]~q ;
wire \cpu|M_alu_result[16]~q ;
wire \cpu|M_alu_result[15]~q ;
wire \cpu|M_alu_result[14]~q ;
wire \cpu|M_alu_result[13]~q ;
wire \mm_interconnect_0|router|Equal1~0_combout ;
wire \cpu|M_alu_result[12]~q ;
wire \cpu|M_alu_result[11]~q ;
wire \cpu|M_alu_result[10]~q ;
wire \cpu|M_alu_result[9]~q ;
wire \cpu|M_alu_result[8]~q ;
wire \cpu|M_alu_result[7]~q ;
wire \mm_interconnect_0|router|Equal2~0_combout ;
wire \mm_interconnect_0|router|Equal4~0_combout ;
wire \mm_interconnect_0|led_pio_s1_translator|wait_latency_counter[1]~q ;
wire \mm_interconnect_0|led_pio_s1_translator|wait_latency_counter[0]~q ;
wire \cpu|M_alu_result[3]~q ;
wire \cpu|M_alu_result[2]~q ;
wire \cpu|M_st_data[1]~q ;
wire \cpu|M_st_data[2]~q ;
wire \cpu|M_st_data[3]~q ;
wire \cpu|M_st_data[4]~q ;
wire \cpu|M_st_data[5]~q ;
wire \cpu|M_st_data[6]~q ;
wire \cpu|M_st_data[7]~q ;
wire \cpu|d_read~q ;
wire \mm_interconnect_0|rsp_mux|WideOr1~combout ;
wire \mm_interconnect_0|cpu_data_master_translator|read_accepted~q ;
wire \mm_interconnect_0|sys_clk_timer_s1_agent_rsp_fifo|mem_used[1]~q ;
wire \mm_interconnect_0|sys_clk_timer_s1_translator|wait_latency_counter[1]~q ;
wire \mm_interconnect_0|sys_clk_timer_s1_translator|wait_latency_counter[0]~q ;
wire \jtag_uart|av_waitrequest~q ;
wire \mm_interconnect_0|router|Equal6~0_combout ;
wire \mm_interconnect_0|cmd_mux_002|saved_grant[0]~q ;
wire \cpu|the_processor_cpu_nios2_oci|the_processor_cpu_nios2_ocimem|waitrequest~q ;
wire \mm_interconnect_0|cpu_jtag_debug_module_agent_rsp_fifo|mem_used[1]~q ;
wire \mm_interconnect_0|cmd_mux_003|saved_grant[0]~q ;
wire \mm_interconnect_0|onchip_mem_s1_agent_rsp_fifo|mem_used[1]~q ;
wire \mm_interconnect_0|cpu_data_master_translator|read_accepted~0_combout ;
wire \cpu|hbreak_enabled~q ;
wire \mm_interconnect_0|cpu_data_master_translator|uav_read~0_combout ;
wire \mm_interconnect_0|cmd_demux|src2_valid~2_combout ;
wire \mm_interconnect_0|cmd_mux_002|saved_grant[1]~q ;
wire \cpu|i_read~q ;
wire \mm_interconnect_0|cpu_instruction_master_limiter|has_pending_responses~q ;
wire \cpu|ic_fill_tag[5]~q ;
wire \cpu|ic_fill_tag[4]~q ;
wire \cpu|ic_fill_tag[3]~q ;
wire \cpu|ic_fill_tag[2]~q ;
wire \cpu|ic_fill_tag[1]~q ;
wire \cpu|ic_fill_tag[0]~q ;
wire \mm_interconnect_0|router_001|Equal1~0_combout ;
wire \mm_interconnect_0|cmd_demux_001|src0_valid~0_combout ;
wire \mm_interconnect_0|cpu_jtag_debug_module_agent|rf_source_valid~0_combout ;
wire \mm_interconnect_0|cmd_demux|src3_valid~0_combout ;
wire \mm_interconnect_0|cmd_mux_003|saved_grant[1]~q ;
wire \mm_interconnect_0|cpu_instruction_master_limiter|last_dest_id[1]~q ;
wire \mm_interconnect_0|cmd_demux_001|src1_valid~0_combout ;
wire \mm_interconnect_0|jtag_uart_avalon_jtag_slave_translator|read_latency_shift_reg~0_combout ;
wire \sys_clk_timer|period_l_wr_strobe~0_combout ;
wire \mm_interconnect_0|rsp_mux|src_data[0]~combout ;
wire \mm_interconnect_0|rsp_mux|src_payload~1_combout ;
wire \mm_interconnect_0|rsp_mux|src_data[8]~combout ;
wire \mm_interconnect_0|rsp_mux|src_payload~2_combout ;
wire \mm_interconnect_0|cmd_demux_001|WideOr0~0_combout ;
wire \mm_interconnect_0|cpu_instruction_master_limiter|nonposted_cmd_accepted~combout ;
wire \cpu|ic_fill_line[5]~q ;
wire \mm_interconnect_0|cmd_mux_002|src_data[46]~combout ;
wire \mm_interconnect_0|rsp_mux|src_data[5]~combout ;
wire \mm_interconnect_0|rsp_mux|src_payload~4_combout ;
wire \mm_interconnect_0|rsp_mux|src_payload~6_combout ;
wire \mm_interconnect_0|rsp_mux|src_payload~7_combout ;
wire \mm_interconnect_0|rsp_mux|src_data[4]~combout ;
wire \mm_interconnect_0|rsp_mux|src_payload~9_combout ;
wire \mm_interconnect_0|rsp_mux|src_payload~11_combout ;
wire \mm_interconnect_0|rsp_mux|src_payload~12_combout ;
wire \mm_interconnect_0|rsp_mux|src_data[6]~combout ;
wire \mm_interconnect_0|rsp_mux|src_payload~14_combout ;
wire \mm_interconnect_0|rsp_mux|src_payload~16_combout ;
wire \mm_interconnect_0|rsp_mux|src_payload~17_combout ;
wire \mm_interconnect_0|rsp_mux|src_data[7]~combout ;
wire \mm_interconnect_0|rsp_mux|src_payload~18_combout ;
wire \mm_interconnect_0|rsp_mux|src_payload~20_combout ;
wire \mm_interconnect_0|rsp_mux|src_payload~21_combout ;
wire \jtag_uart|ien_AE~q ;
wire \jtag_uart|av_readdata[9]~combout ;
wire \jtag_uart|ien_AF~q ;
wire \jtag_uart|av_readdata[8]~0_combout ;
wire \mm_interconnect_0|rsp_mux|src_payload~22_combout ;
wire \mm_interconnect_0|rsp_mux|src_payload~23_combout ;
wire \mm_interconnect_0|rsp_mux|src_payload~25_combout ;
wire \mm_interconnect_0|rsp_mux|src_payload~26_combout ;
wire \mm_interconnect_0|rsp_mux|src_payload~27_combout ;
wire \mm_interconnect_0|rsp_mux|src_data[9]~combout ;
wire \mm_interconnect_0|rsp_mux|src_data[3]~combout ;
wire \mm_interconnect_0|rsp_mux|src_payload~29_combout ;
wire \mm_interconnect_0|rsp_mux|src_data[2]~combout ;
wire \mm_interconnect_0|rsp_mux|src_payload~30_combout ;
wire \mm_interconnect_0|rsp_mux|src_data[1]~combout ;
wire \mm_interconnect_0|rsp_mux|src_payload~32_combout ;
wire \rst_controller|r_early_rst~q ;
wire \jtag_uart|the_processor_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|b_full~q ;
wire \sys_clk_timer|timeout_occurred~q ;
wire \sys_clk_timer|control_register[0]~q ;
wire \cpu|ic_fill_line[0]~q ;
wire \cpu|ic_fill_line[1]~q ;
wire \cpu|ic_fill_line[2]~q ;
wire \cpu|ic_fill_line[3]~q ;
wire \cpu|ic_fill_line[4]~q ;
wire \mm_interconnect_0|cmd_mux_003|src_payload~0_combout ;
wire \cpu|ic_fill_ap_offset[0]~q ;
wire \mm_interconnect_0|cmd_mux_003|src_data[38]~combout ;
wire \cpu|ic_fill_ap_offset[1]~q ;
wire \mm_interconnect_0|cmd_mux_003|src_data[39]~combout ;
wire \cpu|ic_fill_ap_offset[2]~q ;
wire \mm_interconnect_0|cmd_mux_003|src_data[40]~combout ;
wire \mm_interconnect_0|cmd_mux_003|src_data[41]~combout ;
wire \mm_interconnect_0|cmd_mux_003|src_data[42]~combout ;
wire \mm_interconnect_0|cmd_mux_003|src_data[43]~combout ;
wire \mm_interconnect_0|cmd_mux_003|src_data[44]~combout ;
wire \mm_interconnect_0|cmd_mux_003|src_data[45]~combout ;
wire \mm_interconnect_0|cmd_mux_003|src_data[46]~combout ;
wire \mm_interconnect_0|cmd_mux_003|src_data[47]~combout ;
wire \mm_interconnect_0|cmd_mux_003|src_data[48]~combout ;
wire \mm_interconnect_0|cmd_mux_003|src_data[49]~combout ;
wire \mm_interconnect_0|cmd_mux_003|src_data[50]~combout ;
wire \cpu|M_mem_byte_en[0]~q ;
wire \mm_interconnect_0|cmd_mux_003|src_data[32]~combout ;
wire \switches_pio|readdata[0]~q ;
wire \led_pio|readdata[0]~combout ;
wire \jtag_uart|read_0~q ;
wire \sys_clk_timer|readdata[0]~q ;
wire \jtag_uart|the_processor_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[0]~q ;
wire \mm_interconnect_0|cmd_mux_003|src_payload~1_combout ;
wire \cpu|M_mem_byte_en[2]~q ;
wire \mm_interconnect_0|cmd_mux_003|src_data[34]~combout ;
wire \mm_interconnect_0|cmd_mux_003|src_payload~2_combout ;
wire \cpu|M_mem_byte_en[1]~q ;
wire \mm_interconnect_0|cmd_mux_003|src_data[33]~combout ;
wire \led_pio|readdata[8]~combout ;
wire \sys_clk_timer|readdata[8]~q ;
wire \switches_pio|readdata[8]~q ;
wire \cpu|M_st_data[24]~q ;
wire \mm_interconnect_0|cmd_mux_003|src_payload~3_combout ;
wire \cpu|M_mem_byte_en[3]~q ;
wire \mm_interconnect_0|cmd_mux_003|src_data[35]~combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~0_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_data[38]~combout ;
wire \mm_interconnect_0|cmd_mux_002|src_data[41]~combout ;
wire \mm_interconnect_0|cmd_mux_002|src_data[40]~combout ;
wire \mm_interconnect_0|cmd_mux_002|src_data[39]~combout ;
wire \mm_interconnect_0|cmd_mux_002|src_data[45]~combout ;
wire \mm_interconnect_0|cmd_mux_002|src_data[44]~combout ;
wire \mm_interconnect_0|cmd_mux_002|src_data[43]~combout ;
wire \mm_interconnect_0|cmd_mux_002|src_data[42]~combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~1_combout ;
wire \mm_interconnect_0|cmd_mux_003|src_payload~4_combout ;
wire \switches_pio|readdata[5]~q ;
wire \led_pio|readdata[5]~combout ;
wire \sys_clk_timer|readdata[5]~q ;
wire \mm_interconnect_0|cmd_mux_003|src_payload~5_combout ;
wire \jtag_uart|the_processor_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[5]~q ;
wire \mm_interconnect_0|cmd_mux_003|src_payload~6_combout ;
wire \jtag_uart|the_processor_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|b_full~q ;
wire \sys_clk_timer|readdata[13]~q ;
wire \cpu|M_st_data[29]~q ;
wire \mm_interconnect_0|cmd_mux_003|src_payload~7_combout ;
wire \mm_interconnect_0|cmd_mux_003|src_payload~8_combout ;
wire \switches_pio|readdata[4]~q ;
wire \led_pio|readdata[4]~combout ;
wire \sys_clk_timer|readdata[4]~q ;
wire \mm_interconnect_0|cmd_mux_003|src_payload~9_combout ;
wire \jtag_uart|the_processor_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[4]~q ;
wire \mm_interconnect_0|cmd_mux_003|src_payload~10_combout ;
wire \jtag_uart|the_processor_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|b_non_empty~q ;
wire \sys_clk_timer|readdata[12]~q ;
wire \cpu|M_st_data[28]~q ;
wire \mm_interconnect_0|cmd_mux_003|src_payload~11_combout ;
wire \mm_interconnect_0|cmd_mux_003|src_payload~12_combout ;
wire \switches_pio|readdata[6]~q ;
wire \led_pio|readdata[6]~combout ;
wire \sys_clk_timer|readdata[6]~q ;
wire \mm_interconnect_0|cmd_mux_003|src_payload~13_combout ;
wire \mm_interconnect_0|cmd_mux_003|src_payload~14_combout ;
wire \jtag_uart|woverflow~q ;
wire \sys_clk_timer|readdata[14]~q ;
wire \cpu|M_st_data[30]~q ;
wire \mm_interconnect_0|cmd_mux_003|src_payload~15_combout ;
wire \mm_interconnect_0|cmd_mux_003|src_payload~16_combout ;
wire \switches_pio|readdata[7]~q ;
wire \led_pio|readdata[7]~combout ;
wire \sys_clk_timer|readdata[7]~q ;
wire \mm_interconnect_0|cmd_mux_003|src_payload~17_combout ;
wire \mm_interconnect_0|cmd_mux_003|src_payload~18_combout ;
wire \jtag_uart|rvalid~q ;
wire \sys_clk_timer|readdata[15]~q ;
wire \cpu|M_st_data[31]~q ;
wire \mm_interconnect_0|cmd_mux_003|src_payload~19_combout ;
wire \mm_interconnect_0|cmd_mux_003|src_payload~20_combout ;
wire \sys_clk_timer|readdata[11]~q ;
wire \cpu|M_st_data[27]~q ;
wire \mm_interconnect_0|cmd_mux_003|src_payload~21_combout ;
wire \mm_interconnect_0|cmd_mux_003|src_payload~22_combout ;
wire \jtag_uart|ac~q ;
wire \sys_clk_timer|readdata[10]~q ;
wire \cpu|M_st_data[26]~q ;
wire \mm_interconnect_0|cmd_mux_003|src_payload~23_combout ;
wire \cpu|M_st_data[25]~q ;
wire \mm_interconnect_0|cmd_mux_003|src_payload~24_combout ;
wire \mm_interconnect_0|cmd_mux_003|src_payload~25_combout ;
wire \led_pio|readdata[9]~combout ;
wire \sys_clk_timer|readdata[9]~q ;
wire \switches_pio|readdata[9]~q ;
wire \mm_interconnect_0|cmd_mux_003|src_payload~26_combout ;
wire \led_pio|readdata[3]~combout ;
wire \sys_clk_timer|readdata[3]~q ;
wire \switches_pio|readdata[3]~q ;
wire \mm_interconnect_0|cmd_mux_003|src_payload~27_combout ;
wire \jtag_uart|the_processor_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[3]~q ;
wire \mm_interconnect_0|cmd_mux_003|src_payload~28_combout ;
wire \led_pio|readdata[2]~combout ;
wire \sys_clk_timer|readdata[2]~q ;
wire \switches_pio|readdata[2]~q ;
wire \jtag_uart|the_processor_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[2]~q ;
wire \mm_interconnect_0|cmd_mux_003|src_payload~29_combout ;
wire \mm_interconnect_0|cmd_mux_003|src_payload~30_combout ;
wire \led_pio|readdata[1]~combout ;
wire \sys_clk_timer|readdata[1]~q ;
wire \switches_pio|readdata[1]~q ;
wire \mm_interconnect_0|cmd_mux_003|src_payload~31_combout ;
wire \jtag_uart|the_processor_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[1]~q ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~2_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_data[32]~combout ;
wire \mm_interconnect_0|rsp_mux_001|WideOr1~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[24]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[0]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[1]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[2]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[3]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[4]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[5]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[22]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[23]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[25]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[26]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[14]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[12]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[11]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[16]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[15]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[13]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[21]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[29]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[27]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[28]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[30]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[31]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[10]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[6]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[8]~combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~3_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[7]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[20]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[19]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[18]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[17]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[9]~combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~4_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~5_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_data[34]~combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~6_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_data[33]~combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~7_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_data[35]~combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~8_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~9_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~10_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~11_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~12_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~13_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~14_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~15_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~16_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~17_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~18_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~19_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~20_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~21_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~22_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~23_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~24_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~25_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~26_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~27_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~28_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~29_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~30_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~31_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~32_combout ;
wire \rst_controller|alt_rst_req_sync_uq1|altera_reset_synchronizer_int_chain[1]~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_1[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~14_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~6_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~6_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~7_combout ;
wire \auto_hub|~GND~combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~_wirecell_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~_wirecell_combout ;
wire \clk_clk~input_o ;
wire \switches_pio_external_connection_export[0]~input_o ;
wire \switches_pio_external_connection_export[8]~input_o ;
wire \switches_pio_external_connection_export[5]~input_o ;
wire \switches_pio_external_connection_export[4]~input_o ;
wire \switches_pio_external_connection_export[6]~input_o ;
wire \switches_pio_external_connection_export[7]~input_o ;
wire \switches_pio_external_connection_export[9]~input_o ;
wire \switches_pio_external_connection_export[3]~input_o ;
wire \switches_pio_external_connection_export[2]~input_o ;
wire \switches_pio_external_connection_export[1]~input_o ;
wire \reset_reset_n~input_o ;
wire \altera_reserved_tms~input_o ;
wire \altera_reserved_tck~input_o ;
wire \altera_reserved_tdi~input_o ;
wire \altera_internal_jtag~TCKUTAP ;
wire \altera_internal_jtag~TMSUTAP ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~6_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~7_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~9_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~12_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~13_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~10_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~11_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ;
wire \altera_internal_jtag~TDIUTAP ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal1~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ;
wire \~GND~combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~8_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~6_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~7_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal11~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg_proc~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_tdo_sel_reg[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_tdo_sel_reg[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~8_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~6_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~7_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~6_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~8_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~9_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~7_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~6_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~7_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~q ;
wire \altera_internal_jtag~TDO ;


processor_processor_cpu cpu(
	.M_st_data_8(\cpu|M_st_data[8]~q ),
	.M_st_data_9(\cpu|M_st_data[9]~q ),
	.readdata_0(\cpu|the_processor_cpu_nios2_oci|readdata[0]~q ),
	.readdata_16(\cpu|the_processor_cpu_nios2_oci|readdata[16]~q ),
	.M_st_data_16(\cpu|M_st_data[16]~q ),
	.readdata_8(\cpu|the_processor_cpu_nios2_oci|readdata[8]~q ),
	.readdata_24(\cpu|the_processor_cpu_nios2_oci|readdata[24]~q ),
	.readdata_5(\cpu|the_processor_cpu_nios2_oci|readdata[5]~q ),
	.readdata_21(\cpu|the_processor_cpu_nios2_oci|readdata[21]~q ),
	.M_st_data_21(\cpu|M_st_data[21]~q ),
	.readdata_13(\cpu|the_processor_cpu_nios2_oci|readdata[13]~q ),
	.M_st_data_13(\cpu|M_st_data[13]~q ),
	.readdata_29(\cpu|the_processor_cpu_nios2_oci|readdata[29]~q ),
	.readdata_4(\cpu|the_processor_cpu_nios2_oci|readdata[4]~q ),
	.readdata_20(\cpu|the_processor_cpu_nios2_oci|readdata[20]~q ),
	.M_st_data_20(\cpu|M_st_data[20]~q ),
	.readdata_12(\cpu|the_processor_cpu_nios2_oci|readdata[12]~q ),
	.M_st_data_12(\cpu|M_st_data[12]~q ),
	.readdata_28(\cpu|the_processor_cpu_nios2_oci|readdata[28]~q ),
	.readdata_6(\cpu|the_processor_cpu_nios2_oci|readdata[6]~q ),
	.readdata_22(\cpu|the_processor_cpu_nios2_oci|readdata[22]~q ),
	.M_st_data_22(\cpu|M_st_data[22]~q ),
	.readdata_14(\cpu|the_processor_cpu_nios2_oci|readdata[14]~q ),
	.M_st_data_14(\cpu|M_st_data[14]~q ),
	.readdata_30(\cpu|the_processor_cpu_nios2_oci|readdata[30]~q ),
	.readdata_7(\cpu|the_processor_cpu_nios2_oci|readdata[7]~q ),
	.readdata_23(\cpu|the_processor_cpu_nios2_oci|readdata[23]~q ),
	.M_st_data_23(\cpu|M_st_data[23]~q ),
	.readdata_15(\cpu|the_processor_cpu_nios2_oci|readdata[15]~q ),
	.M_st_data_15(\cpu|M_st_data[15]~q ),
	.readdata_31(\cpu|the_processor_cpu_nios2_oci|readdata[31]~q ),
	.readdata_11(\cpu|the_processor_cpu_nios2_oci|readdata[11]~q ),
	.M_st_data_11(\cpu|M_st_data[11]~q ),
	.readdata_27(\cpu|the_processor_cpu_nios2_oci|readdata[27]~q ),
	.readdata_10(\cpu|the_processor_cpu_nios2_oci|readdata[10]~q ),
	.M_st_data_10(\cpu|M_st_data[10]~q ),
	.readdata_26(\cpu|the_processor_cpu_nios2_oci|readdata[26]~q ),
	.readdata_25(\cpu|the_processor_cpu_nios2_oci|readdata[25]~q ),
	.readdata_9(\cpu|the_processor_cpu_nios2_oci|readdata[9]~q ),
	.readdata_3(\cpu|the_processor_cpu_nios2_oci|readdata[3]~q ),
	.readdata_19(\cpu|the_processor_cpu_nios2_oci|readdata[19]~q ),
	.M_st_data_19(\cpu|M_st_data[19]~q ),
	.readdata_2(\cpu|the_processor_cpu_nios2_oci|readdata[2]~q ),
	.readdata_18(\cpu|the_processor_cpu_nios2_oci|readdata[18]~q ),
	.M_st_data_18(\cpu|M_st_data[18]~q ),
	.readdata_1(\cpu|the_processor_cpu_nios2_oci|readdata[1]~q ),
	.readdata_17(\cpu|the_processor_cpu_nios2_oci|readdata[17]~q ),
	.M_st_data_17(\cpu|M_st_data[17]~q ),
	.sr_0(\cpu|the_processor_cpu_nios2_oci|the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_tck|sr[0]~q ),
	.ir_out_0(\cpu|the_processor_cpu_nios2_oci|the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_tck|ir_out[0]~q ),
	.ir_out_1(\cpu|the_processor_cpu_nios2_oci|the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_tck|ir_out[1]~q ),
	.M_st_data_0(\cpu|M_st_data[0]~q ),
	.r_sync_rst(\rst_controller|r_sync_rst~q ),
	.clr_break_line1(\cpu|clr_break_line~q ),
	.d_write1(\cpu|d_write~q ),
	.M_alu_result_5(\cpu|M_alu_result[5]~q ),
	.M_alu_result_4(\cpu|M_alu_result[4]~q ),
	.M_alu_result_6(\cpu|M_alu_result[6]~q ),
	.M_alu_result_16(\cpu|M_alu_result[16]~q ),
	.M_alu_result_15(\cpu|M_alu_result[15]~q ),
	.M_alu_result_14(\cpu|M_alu_result[14]~q ),
	.M_alu_result_13(\cpu|M_alu_result[13]~q ),
	.M_alu_result_12(\cpu|M_alu_result[12]~q ),
	.M_alu_result_11(\cpu|M_alu_result[11]~q ),
	.M_alu_result_10(\cpu|M_alu_result[10]~q ),
	.M_alu_result_9(\cpu|M_alu_result[9]~q ),
	.M_alu_result_8(\cpu|M_alu_result[8]~q ),
	.M_alu_result_7(\cpu|M_alu_result[7]~q ),
	.M_alu_result_3(\cpu|M_alu_result[3]~q ),
	.M_alu_result_2(\cpu|M_alu_result[2]~q ),
	.M_st_data_1(\cpu|M_st_data[1]~q ),
	.M_st_data_2(\cpu|M_st_data[2]~q ),
	.M_st_data_3(\cpu|M_st_data[3]~q ),
	.M_st_data_4(\cpu|M_st_data[4]~q ),
	.M_st_data_5(\cpu|M_st_data[5]~q ),
	.M_st_data_6(\cpu|M_st_data[6]~q ),
	.M_st_data_7(\cpu|M_st_data[7]~q ),
	.d_read1(\cpu|d_read~q ),
	.WideOr1(\mm_interconnect_0|rsp_mux|WideOr1~combout ),
	.saved_grant_0(\mm_interconnect_0|cmd_mux_002|saved_grant[0]~q ),
	.jtag_debug_module_waitrequest(\cpu|the_processor_cpu_nios2_oci|the_processor_cpu_nios2_ocimem|waitrequest~q ),
	.mem_used_1(\mm_interconnect_0|cpu_jtag_debug_module_agent_rsp_fifo|mem_used[1]~q ),
	.read_accepted(\mm_interconnect_0|cpu_data_master_translator|read_accepted~0_combout ),
	.hbreak_enabled1(\cpu|hbreak_enabled~q ),
	.src2_valid(\mm_interconnect_0|cmd_demux|src2_valid~2_combout ),
	.saved_grant_1(\mm_interconnect_0|cmd_mux_002|saved_grant[1]~q ),
	.i_read1(\cpu|i_read~q ),
	.has_pending_responses(\mm_interconnect_0|cpu_instruction_master_limiter|has_pending_responses~q ),
	.ic_fill_tag_5(\cpu|ic_fill_tag[5]~q ),
	.ic_fill_tag_4(\cpu|ic_fill_tag[4]~q ),
	.ic_fill_tag_3(\cpu|ic_fill_tag[3]~q ),
	.ic_fill_tag_2(\cpu|ic_fill_tag[2]~q ),
	.ic_fill_tag_1(\cpu|ic_fill_tag[1]~q ),
	.ic_fill_tag_0(\cpu|ic_fill_tag[0]~q ),
	.Equal1(\mm_interconnect_0|router_001|Equal1~0_combout ),
	.src0_valid(\mm_interconnect_0|cmd_demux_001|src0_valid~0_combout ),
	.rf_source_valid(\mm_interconnect_0|cpu_jtag_debug_module_agent|rf_source_valid~0_combout ),
	.last_dest_id_1(\mm_interconnect_0|cpu_instruction_master_limiter|last_dest_id[1]~q ),
	.d_readdata({\mm_interconnect_0|rsp_mux|src_payload~21_combout ,\mm_interconnect_0|rsp_mux|src_payload~17_combout ,\mm_interconnect_0|rsp_mux|src_payload~7_combout ,\mm_interconnect_0|rsp_mux|src_payload~12_combout ,\mm_interconnect_0|rsp_mux|src_payload~23_combout ,
\mm_interconnect_0|rsp_mux|src_payload~26_combout ,\mm_interconnect_0|rsp_mux|src_payload~27_combout ,\mm_interconnect_0|rsp_mux|src_payload~2_combout ,\mm_interconnect_0|rsp_mux|src_payload~18_combout ,\mm_interconnect_0|rsp_mux|src_payload~14_combout ,
\mm_interconnect_0|rsp_mux|src_payload~4_combout ,\mm_interconnect_0|rsp_mux|src_payload~9_combout ,\mm_interconnect_0|rsp_mux|src_payload~29_combout ,\mm_interconnect_0|rsp_mux|src_payload~30_combout ,\mm_interconnect_0|rsp_mux|src_payload~32_combout ,
\mm_interconnect_0|rsp_mux|src_payload~1_combout ,\mm_interconnect_0|rsp_mux|src_payload~20_combout ,\mm_interconnect_0|rsp_mux|src_payload~16_combout ,\mm_interconnect_0|rsp_mux|src_payload~6_combout ,\mm_interconnect_0|rsp_mux|src_payload~11_combout ,
\mm_interconnect_0|rsp_mux|src_payload~22_combout ,\mm_interconnect_0|rsp_mux|src_payload~25_combout ,\mm_interconnect_0|rsp_mux|src_data[9]~combout ,\mm_interconnect_0|rsp_mux|src_data[8]~combout ,\mm_interconnect_0|rsp_mux|src_data[7]~combout ,
\mm_interconnect_0|rsp_mux|src_data[6]~combout ,\mm_interconnect_0|rsp_mux|src_data[5]~combout ,\mm_interconnect_0|rsp_mux|src_data[4]~combout ,\mm_interconnect_0|rsp_mux|src_data[3]~combout ,\mm_interconnect_0|rsp_mux|src_data[2]~combout ,
\mm_interconnect_0|rsp_mux|src_data[1]~combout ,\mm_interconnect_0|rsp_mux|src_data[0]~combout }),
	.WideOr0(\mm_interconnect_0|cmd_demux_001|WideOr0~0_combout ),
	.nonposted_cmd_accepted(\mm_interconnect_0|cpu_instruction_master_limiter|nonposted_cmd_accepted~combout ),
	.ic_fill_line_5(\cpu|ic_fill_line[5]~q ),
	.src_data_46(\mm_interconnect_0|cmd_mux_002|src_data[46]~combout ),
	.av_readdata_9(\jtag_uart|av_readdata[9]~combout ),
	.av_readdata_8(\jtag_uart|av_readdata[8]~0_combout ),
	.r_early_rst(\rst_controller|r_early_rst~q ),
	.timeout_occurred(\sys_clk_timer|timeout_occurred~q ),
	.control_register_0(\sys_clk_timer|control_register[0]~q ),
	.ic_fill_line_0(\cpu|ic_fill_line[0]~q ),
	.ic_fill_line_1(\cpu|ic_fill_line[1]~q ),
	.ic_fill_line_2(\cpu|ic_fill_line[2]~q ),
	.ic_fill_line_3(\cpu|ic_fill_line[3]~q ),
	.ic_fill_line_4(\cpu|ic_fill_line[4]~q ),
	.ic_fill_ap_offset_0(\cpu|ic_fill_ap_offset[0]~q ),
	.ic_fill_ap_offset_1(\cpu|ic_fill_ap_offset[1]~q ),
	.ic_fill_ap_offset_2(\cpu|ic_fill_ap_offset[2]~q ),
	.M_mem_byte_en_0(\cpu|M_mem_byte_en[0]~q ),
	.M_mem_byte_en_2(\cpu|M_mem_byte_en[2]~q ),
	.M_mem_byte_en_1(\cpu|M_mem_byte_en[1]~q ),
	.M_st_data_24(\cpu|M_st_data[24]~q ),
	.M_mem_byte_en_3(\cpu|M_mem_byte_en[3]~q ),
	.src_payload(\mm_interconnect_0|cmd_mux_002|src_payload~0_combout ),
	.src_data_38(\mm_interconnect_0|cmd_mux_002|src_data[38]~combout ),
	.src_data_41(\mm_interconnect_0|cmd_mux_002|src_data[41]~combout ),
	.src_data_40(\mm_interconnect_0|cmd_mux_002|src_data[40]~combout ),
	.src_data_39(\mm_interconnect_0|cmd_mux_002|src_data[39]~combout ),
	.src_data_45(\mm_interconnect_0|cmd_mux_002|src_data[45]~combout ),
	.src_data_44(\mm_interconnect_0|cmd_mux_002|src_data[44]~combout ),
	.src_data_43(\mm_interconnect_0|cmd_mux_002|src_data[43]~combout ),
	.src_data_42(\mm_interconnect_0|cmd_mux_002|src_data[42]~combout ),
	.src_payload1(\mm_interconnect_0|cmd_mux_002|src_payload~1_combout ),
	.M_st_data_29(\cpu|M_st_data[29]~q ),
	.M_st_data_28(\cpu|M_st_data[28]~q ),
	.M_st_data_30(\cpu|M_st_data[30]~q ),
	.M_st_data_31(\cpu|M_st_data[31]~q ),
	.M_st_data_27(\cpu|M_st_data[27]~q ),
	.M_st_data_26(\cpu|M_st_data[26]~q ),
	.M_st_data_25(\cpu|M_st_data[25]~q ),
	.src_payload2(\mm_interconnect_0|cmd_mux_002|src_payload~2_combout ),
	.src_data_32(\mm_interconnect_0|cmd_mux_002|src_data[32]~combout ),
	.WideOr11(\mm_interconnect_0|rsp_mux_001|WideOr1~combout ),
	.i_readdata({\mm_interconnect_0|rsp_mux_001|src_data[31]~combout ,\mm_interconnect_0|rsp_mux_001|src_data[30]~combout ,\mm_interconnect_0|rsp_mux_001|src_data[29]~combout ,\mm_interconnect_0|rsp_mux_001|src_data[28]~combout ,
\mm_interconnect_0|rsp_mux_001|src_data[27]~combout ,\mm_interconnect_0|rsp_mux_001|src_data[26]~combout ,\mm_interconnect_0|rsp_mux_001|src_data[25]~combout ,\mm_interconnect_0|rsp_mux_001|src_data[24]~combout ,
\mm_interconnect_0|rsp_mux_001|src_data[23]~combout ,\mm_interconnect_0|rsp_mux_001|src_data[22]~combout ,\mm_interconnect_0|rsp_mux_001|src_data[21]~combout ,\mm_interconnect_0|rsp_mux_001|src_data[20]~combout ,
\mm_interconnect_0|rsp_mux_001|src_data[19]~combout ,\mm_interconnect_0|rsp_mux_001|src_data[18]~combout ,\mm_interconnect_0|rsp_mux_001|src_data[17]~combout ,\mm_interconnect_0|rsp_mux_001|src_data[16]~combout ,
\mm_interconnect_0|rsp_mux_001|src_data[15]~combout ,\mm_interconnect_0|rsp_mux_001|src_data[14]~combout ,\mm_interconnect_0|rsp_mux_001|src_data[13]~combout ,\mm_interconnect_0|rsp_mux_001|src_data[12]~combout ,
\mm_interconnect_0|rsp_mux_001|src_data[11]~combout ,\mm_interconnect_0|rsp_mux_001|src_data[10]~combout ,\mm_interconnect_0|rsp_mux_001|src_data[9]~combout ,\mm_interconnect_0|rsp_mux_001|src_data[8]~combout ,
\mm_interconnect_0|rsp_mux_001|src_data[7]~combout ,\mm_interconnect_0|rsp_mux_001|src_data[6]~combout ,\mm_interconnect_0|rsp_mux_001|src_data[5]~combout ,\mm_interconnect_0|rsp_mux_001|src_data[4]~combout ,\mm_interconnect_0|rsp_mux_001|src_data[3]~combout ,
\mm_interconnect_0|rsp_mux_001|src_data[2]~combout ,\mm_interconnect_0|rsp_mux_001|src_data[1]~combout ,\mm_interconnect_0|rsp_mux_001|src_data[0]~combout }),
	.src_payload3(\mm_interconnect_0|cmd_mux_002|src_payload~3_combout ),
	.src_payload4(\mm_interconnect_0|cmd_mux_002|src_payload~4_combout ),
	.src_payload5(\mm_interconnect_0|cmd_mux_002|src_payload~5_combout ),
	.src_data_34(\mm_interconnect_0|cmd_mux_002|src_data[34]~combout ),
	.src_payload6(\mm_interconnect_0|cmd_mux_002|src_payload~6_combout ),
	.src_data_33(\mm_interconnect_0|cmd_mux_002|src_data[33]~combout ),
	.src_payload7(\mm_interconnect_0|cmd_mux_002|src_payload~7_combout ),
	.src_data_35(\mm_interconnect_0|cmd_mux_002|src_data[35]~combout ),
	.src_payload8(\mm_interconnect_0|cmd_mux_002|src_payload~8_combout ),
	.src_payload9(\mm_interconnect_0|cmd_mux_002|src_payload~9_combout ),
	.src_payload10(\mm_interconnect_0|cmd_mux_002|src_payload~10_combout ),
	.src_payload11(\mm_interconnect_0|cmd_mux_002|src_payload~11_combout ),
	.src_payload12(\mm_interconnect_0|cmd_mux_002|src_payload~12_combout ),
	.src_payload13(\mm_interconnect_0|cmd_mux_002|src_payload~13_combout ),
	.src_payload14(\mm_interconnect_0|cmd_mux_002|src_payload~14_combout ),
	.src_payload15(\mm_interconnect_0|cmd_mux_002|src_payload~15_combout ),
	.src_payload16(\mm_interconnect_0|cmd_mux_002|src_payload~16_combout ),
	.src_payload17(\mm_interconnect_0|cmd_mux_002|src_payload~17_combout ),
	.src_payload18(\mm_interconnect_0|cmd_mux_002|src_payload~18_combout ),
	.src_payload19(\mm_interconnect_0|cmd_mux_002|src_payload~19_combout ),
	.src_payload20(\mm_interconnect_0|cmd_mux_002|src_payload~20_combout ),
	.src_payload21(\mm_interconnect_0|cmd_mux_002|src_payload~21_combout ),
	.src_payload22(\mm_interconnect_0|cmd_mux_002|src_payload~22_combout ),
	.src_payload23(\mm_interconnect_0|cmd_mux_002|src_payload~23_combout ),
	.src_payload24(\mm_interconnect_0|cmd_mux_002|src_payload~24_combout ),
	.src_payload25(\mm_interconnect_0|cmd_mux_002|src_payload~25_combout ),
	.src_payload26(\mm_interconnect_0|cmd_mux_002|src_payload~26_combout ),
	.src_payload27(\mm_interconnect_0|cmd_mux_002|src_payload~27_combout ),
	.src_payload28(\mm_interconnect_0|cmd_mux_002|src_payload~28_combout ),
	.src_payload29(\mm_interconnect_0|cmd_mux_002|src_payload~29_combout ),
	.src_payload30(\mm_interconnect_0|cmd_mux_002|src_payload~30_combout ),
	.src_payload31(\mm_interconnect_0|cmd_mux_002|src_payload~31_combout ),
	.src_payload32(\mm_interconnect_0|cmd_mux_002|src_payload~32_combout ),
	.altera_internal_jtag(\altera_internal_jtag~TCKUTAP ),
	.altera_internal_jtag1(\altera_internal_jtag~TDIUTAP ),
	.state_1(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1]~q ),
	.state_4(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.virtual_ir_scan_reg(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.state_3(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.state_8(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.splitter_nodes_receive_1_3(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_1[3]~q ),
	.irf_reg_0_2(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~q ),
	.irf_reg_1_2(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][1]~q ),
	.clk_clk(\clk_clk~input_o ));

processor_processor_jtag_uart jtag_uart(
	.q_b_0(\jtag_uart|the_processor_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[0] ),
	.Add1(\jtag_uart|Add1~1_sumout ),
	.q_b_5(\jtag_uart|the_processor_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[5] ),
	.Add11(\jtag_uart|Add1~5_sumout ),
	.q_b_4(\jtag_uart|the_processor_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[4] ),
	.Add12(\jtag_uart|Add1~9_sumout ),
	.q_b_6(\jtag_uart|the_processor_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[6] ),
	.Add13(\jtag_uart|Add1~13_sumout ),
	.q_b_7(\jtag_uart|the_processor_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[7] ),
	.M_st_data_10(\cpu|M_st_data[10]~q ),
	.q_b_3(\jtag_uart|the_processor_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[3] ),
	.Add14(\jtag_uart|Add1~17_sumout ),
	.q_b_2(\jtag_uart|the_processor_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[2] ),
	.Add15(\jtag_uart|Add1~21_sumout ),
	.q_b_1(\jtag_uart|the_processor_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[1] ),
	.Add16(\jtag_uart|Add1~25_sumout ),
	.tdo(\jtag_uart|processor_jtag_uart_alt_jtag_atlantic|tdo~q ),
	.M_st_data_0(\cpu|M_st_data[0]~q ),
	.r_sync_rst(\rst_controller|r_sync_rst~q ),
	.clr_break_line(\cpu|clr_break_line~q ),
	.d_write(\cpu|d_write~q ),
	.Equal1(\mm_interconnect_0|router|Equal1~0_combout ),
	.Equal2(\mm_interconnect_0|router|Equal2~0_combout ),
	.M_alu_result_2(\cpu|M_alu_result[2]~q ),
	.M_st_data_1(\cpu|M_st_data[1]~q ),
	.M_st_data_2(\cpu|M_st_data[2]~q ),
	.M_st_data_3(\cpu|M_st_data[3]~q ),
	.M_st_data_4(\cpu|M_st_data[4]~q ),
	.M_st_data_5(\cpu|M_st_data[5]~q ),
	.M_st_data_6(\cpu|M_st_data[6]~q ),
	.M_st_data_7(\cpu|M_st_data[7]~q ),
	.d_read(\cpu|d_read~q ),
	.read_accepted(\mm_interconnect_0|cpu_data_master_translator|read_accepted~q ),
	.av_waitrequest1(\jtag_uart|av_waitrequest~q ),
	.Equal6(\mm_interconnect_0|router|Equal6~0_combout ),
	.uav_read(\mm_interconnect_0|cpu_data_master_translator|uav_read~0_combout ),
	.read_latency_shift_reg(\mm_interconnect_0|jtag_uart_avalon_jtag_slave_translator|read_latency_shift_reg~0_combout ),
	.ien_AE1(\jtag_uart|ien_AE~q ),
	.av_readdata_9(\jtag_uart|av_readdata[9]~combout ),
	.ien_AF1(\jtag_uart|ien_AF~q ),
	.av_readdata_8(\jtag_uart|av_readdata[8]~0_combout ),
	.b_full(\jtag_uart|the_processor_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|b_full~q ),
	.read_01(\jtag_uart|read_0~q ),
	.counter_reg_bit_0(\jtag_uart|the_processor_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[0]~q ),
	.counter_reg_bit_5(\jtag_uart|the_processor_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[5]~q ),
	.b_full1(\jtag_uart|the_processor_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|b_full~q ),
	.counter_reg_bit_4(\jtag_uart|the_processor_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[4]~q ),
	.b_non_empty(\jtag_uart|the_processor_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|b_non_empty~q ),
	.woverflow1(\jtag_uart|woverflow~q ),
	.rvalid1(\jtag_uart|rvalid~q ),
	.ac1(\jtag_uart|ac~q ),
	.counter_reg_bit_3(\jtag_uart|the_processor_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[3]~q ),
	.counter_reg_bit_2(\jtag_uart|the_processor_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[2]~q ),
	.counter_reg_bit_1(\jtag_uart|the_processor_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[1]~q ),
	.altera_internal_jtag(\altera_internal_jtag~TCKUTAP ),
	.altera_internal_jtag1(\altera_internal_jtag~TDIUTAP ),
	.state_4(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.splitter_nodes_receive_0_3(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3]~q ),
	.virtual_ir_scan_reg(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.clr_reg(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.state_3(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.state_8(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.irf_reg_0_1(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~q ),
	.clk_clk(\clk_clk~input_o ));

processor_processor_sys_clk_timer sys_clk_timer(
	.writedata({\cpu|M_st_data[15]~q ,\cpu|M_st_data[14]~q ,\cpu|M_st_data[13]~q ,\cpu|M_st_data[12]~q ,\cpu|M_st_data[11]~q ,\cpu|M_st_data[10]~q ,\cpu|M_st_data[9]~q ,\cpu|M_st_data[8]~q ,\cpu|M_st_data[7]~q ,\cpu|M_st_data[6]~q ,\cpu|M_st_data[5]~q ,\cpu|M_st_data[4]~q ,
\cpu|M_st_data[3]~q ,\cpu|M_st_data[2]~q ,\cpu|M_st_data[1]~q ,\cpu|M_st_data[0]~q }),
	.reset_n(\rst_controller|r_sync_rst~q ),
	.clr_break_line(\cpu|clr_break_line~q ),
	.d_write(\cpu|d_write~q ),
	.M_alu_result_5(\cpu|M_alu_result[5]~q ),
	.M_alu_result_4(\cpu|M_alu_result[4]~q ),
	.M_alu_result_6(\cpu|M_alu_result[6]~q ),
	.Equal1(\mm_interconnect_0|router|Equal1~0_combout ),
	.Equal2(\mm_interconnect_0|router|Equal2~0_combout ),
	.M_alu_result_3(\cpu|M_alu_result[3]~q ),
	.M_alu_result_2(\cpu|M_alu_result[2]~q ),
	.mem_used_1(\mm_interconnect_0|sys_clk_timer_s1_agent_rsp_fifo|mem_used[1]~q ),
	.wait_latency_counter_1(\mm_interconnect_0|sys_clk_timer_s1_translator|wait_latency_counter[1]~q ),
	.wait_latency_counter_0(\mm_interconnect_0|sys_clk_timer_s1_translator|wait_latency_counter[0]~q ),
	.period_l_wr_strobe1(\sys_clk_timer|period_l_wr_strobe~0_combout ),
	.timeout_occurred1(\sys_clk_timer|timeout_occurred~q ),
	.control_register_0(\sys_clk_timer|control_register[0]~q ),
	.readdata_0(\sys_clk_timer|readdata[0]~q ),
	.readdata_8(\sys_clk_timer|readdata[8]~q ),
	.readdata_5(\sys_clk_timer|readdata[5]~q ),
	.readdata_13(\sys_clk_timer|readdata[13]~q ),
	.readdata_4(\sys_clk_timer|readdata[4]~q ),
	.readdata_12(\sys_clk_timer|readdata[12]~q ),
	.readdata_6(\sys_clk_timer|readdata[6]~q ),
	.readdata_14(\sys_clk_timer|readdata[14]~q ),
	.readdata_7(\sys_clk_timer|readdata[7]~q ),
	.readdata_15(\sys_clk_timer|readdata[15]~q ),
	.readdata_11(\sys_clk_timer|readdata[11]~q ),
	.readdata_10(\sys_clk_timer|readdata[10]~q ),
	.readdata_9(\sys_clk_timer|readdata[9]~q ),
	.readdata_3(\sys_clk_timer|readdata[3]~q ),
	.readdata_2(\sys_clk_timer|readdata[2]~q ),
	.readdata_1(\sys_clk_timer|readdata[1]~q ),
	.clk(\clk_clk~input_o ));

processor_processor_switches_pio switches_pio(
	.r_sync_rst(\rst_controller|r_sync_rst~q ),
	.M_alu_result_3(\cpu|M_alu_result[3]~q ),
	.M_alu_result_2(\cpu|M_alu_result[2]~q ),
	.readdata_0(\switches_pio|readdata[0]~q ),
	.readdata_8(\switches_pio|readdata[8]~q ),
	.readdata_5(\switches_pio|readdata[5]~q ),
	.readdata_4(\switches_pio|readdata[4]~q ),
	.readdata_6(\switches_pio|readdata[6]~q ),
	.readdata_7(\switches_pio|readdata[7]~q ),
	.readdata_9(\switches_pio|readdata[9]~q ),
	.readdata_3(\switches_pio|readdata[3]~q ),
	.readdata_2(\switches_pio|readdata[2]~q ),
	.readdata_1(\switches_pio|readdata[1]~q ),
	.clk_clk(\clk_clk~input_o ),
	.switches_pio_external_connection_export_0(\switches_pio_external_connection_export[0]~input_o ),
	.switches_pio_external_connection_export_8(\switches_pio_external_connection_export[8]~input_o ),
	.switches_pio_external_connection_export_5(\switches_pio_external_connection_export[5]~input_o ),
	.switches_pio_external_connection_export_4(\switches_pio_external_connection_export[4]~input_o ),
	.switches_pio_external_connection_export_6(\switches_pio_external_connection_export[6]~input_o ),
	.switches_pio_external_connection_export_7(\switches_pio_external_connection_export[7]~input_o ),
	.switches_pio_external_connection_export_9(\switches_pio_external_connection_export[9]~input_o ),
	.switches_pio_external_connection_export_3(\switches_pio_external_connection_export[3]~input_o ),
	.switches_pio_external_connection_export_2(\switches_pio_external_connection_export[2]~input_o ),
	.switches_pio_external_connection_export_1(\switches_pio_external_connection_export[1]~input_o ));

processor_processor_onchip_mem onchip_mem(
	.q_a_0(\onchip_mem|the_altsyncram|auto_generated|q_a[0] ),
	.q_a_16(\onchip_mem|the_altsyncram|auto_generated|q_a[16] ),
	.q_a_8(\onchip_mem|the_altsyncram|auto_generated|q_a[8] ),
	.q_a_24(\onchip_mem|the_altsyncram|auto_generated|q_a[24] ),
	.q_a_5(\onchip_mem|the_altsyncram|auto_generated|q_a[5] ),
	.q_a_21(\onchip_mem|the_altsyncram|auto_generated|q_a[21] ),
	.q_a_13(\onchip_mem|the_altsyncram|auto_generated|q_a[13] ),
	.q_a_29(\onchip_mem|the_altsyncram|auto_generated|q_a[29] ),
	.q_a_4(\onchip_mem|the_altsyncram|auto_generated|q_a[4] ),
	.q_a_20(\onchip_mem|the_altsyncram|auto_generated|q_a[20] ),
	.q_a_12(\onchip_mem|the_altsyncram|auto_generated|q_a[12] ),
	.q_a_28(\onchip_mem|the_altsyncram|auto_generated|q_a[28] ),
	.q_a_6(\onchip_mem|the_altsyncram|auto_generated|q_a[6] ),
	.q_a_22(\onchip_mem|the_altsyncram|auto_generated|q_a[22] ),
	.q_a_14(\onchip_mem|the_altsyncram|auto_generated|q_a[14] ),
	.q_a_30(\onchip_mem|the_altsyncram|auto_generated|q_a[30] ),
	.q_a_7(\onchip_mem|the_altsyncram|auto_generated|q_a[7] ),
	.q_a_23(\onchip_mem|the_altsyncram|auto_generated|q_a[23] ),
	.q_a_15(\onchip_mem|the_altsyncram|auto_generated|q_a[15] ),
	.q_a_31(\onchip_mem|the_altsyncram|auto_generated|q_a[31] ),
	.q_a_11(\onchip_mem|the_altsyncram|auto_generated|q_a[11] ),
	.q_a_27(\onchip_mem|the_altsyncram|auto_generated|q_a[27] ),
	.q_a_10(\onchip_mem|the_altsyncram|auto_generated|q_a[10] ),
	.q_a_26(\onchip_mem|the_altsyncram|auto_generated|q_a[26] ),
	.q_a_25(\onchip_mem|the_altsyncram|auto_generated|q_a[25] ),
	.q_a_9(\onchip_mem|the_altsyncram|auto_generated|q_a[9] ),
	.q_a_3(\onchip_mem|the_altsyncram|auto_generated|q_a[3] ),
	.q_a_19(\onchip_mem|the_altsyncram|auto_generated|q_a[19] ),
	.q_a_2(\onchip_mem|the_altsyncram|auto_generated|q_a[2] ),
	.q_a_18(\onchip_mem|the_altsyncram|auto_generated|q_a[18] ),
	.q_a_1(\onchip_mem|the_altsyncram|auto_generated|q_a[1] ),
	.q_a_17(\onchip_mem|the_altsyncram|auto_generated|q_a[17] ),
	.d_write(\cpu|d_write~q ),
	.saved_grant_0(\mm_interconnect_0|cmd_mux_003|saved_grant[0]~q ),
	.mem_used_1(\mm_interconnect_0|onchip_mem_s1_agent_rsp_fifo|mem_used[1]~q ),
	.src3_valid(\mm_interconnect_0|cmd_demux|src3_valid~0_combout ),
	.saved_grant_1(\mm_interconnect_0|cmd_mux_003|saved_grant[1]~q ),
	.src1_valid(\mm_interconnect_0|cmd_demux_001|src1_valid~0_combout ),
	.r_early_rst(\rst_controller|r_early_rst~q ),
	.src_payload(\mm_interconnect_0|cmd_mux_003|src_payload~0_combout ),
	.src_data_38(\mm_interconnect_0|cmd_mux_003|src_data[38]~combout ),
	.src_data_39(\mm_interconnect_0|cmd_mux_003|src_data[39]~combout ),
	.src_data_40(\mm_interconnect_0|cmd_mux_003|src_data[40]~combout ),
	.src_data_41(\mm_interconnect_0|cmd_mux_003|src_data[41]~combout ),
	.src_data_42(\mm_interconnect_0|cmd_mux_003|src_data[42]~combout ),
	.src_data_43(\mm_interconnect_0|cmd_mux_003|src_data[43]~combout ),
	.src_data_44(\mm_interconnect_0|cmd_mux_003|src_data[44]~combout ),
	.src_data_45(\mm_interconnect_0|cmd_mux_003|src_data[45]~combout ),
	.src_data_46(\mm_interconnect_0|cmd_mux_003|src_data[46]~combout ),
	.src_data_47(\mm_interconnect_0|cmd_mux_003|src_data[47]~combout ),
	.src_data_48(\mm_interconnect_0|cmd_mux_003|src_data[48]~combout ),
	.src_data_49(\mm_interconnect_0|cmd_mux_003|src_data[49]~combout ),
	.src_data_50(\mm_interconnect_0|cmd_mux_003|src_data[50]~combout ),
	.src_data_32(\mm_interconnect_0|cmd_mux_003|src_data[32]~combout ),
	.src_payload1(\mm_interconnect_0|cmd_mux_003|src_payload~1_combout ),
	.src_data_34(\mm_interconnect_0|cmd_mux_003|src_data[34]~combout ),
	.src_payload2(\mm_interconnect_0|cmd_mux_003|src_payload~2_combout ),
	.src_data_33(\mm_interconnect_0|cmd_mux_003|src_data[33]~combout ),
	.src_payload3(\mm_interconnect_0|cmd_mux_003|src_payload~3_combout ),
	.src_data_35(\mm_interconnect_0|cmd_mux_003|src_data[35]~combout ),
	.src_payload4(\mm_interconnect_0|cmd_mux_003|src_payload~4_combout ),
	.src_payload5(\mm_interconnect_0|cmd_mux_003|src_payload~5_combout ),
	.src_payload6(\mm_interconnect_0|cmd_mux_003|src_payload~6_combout ),
	.src_payload7(\mm_interconnect_0|cmd_mux_003|src_payload~7_combout ),
	.src_payload8(\mm_interconnect_0|cmd_mux_003|src_payload~8_combout ),
	.src_payload9(\mm_interconnect_0|cmd_mux_003|src_payload~9_combout ),
	.src_payload10(\mm_interconnect_0|cmd_mux_003|src_payload~10_combout ),
	.src_payload11(\mm_interconnect_0|cmd_mux_003|src_payload~11_combout ),
	.src_payload12(\mm_interconnect_0|cmd_mux_003|src_payload~12_combout ),
	.src_payload13(\mm_interconnect_0|cmd_mux_003|src_payload~13_combout ),
	.src_payload14(\mm_interconnect_0|cmd_mux_003|src_payload~14_combout ),
	.src_payload15(\mm_interconnect_0|cmd_mux_003|src_payload~15_combout ),
	.src_payload16(\mm_interconnect_0|cmd_mux_003|src_payload~16_combout ),
	.src_payload17(\mm_interconnect_0|cmd_mux_003|src_payload~17_combout ),
	.src_payload18(\mm_interconnect_0|cmd_mux_003|src_payload~18_combout ),
	.src_payload19(\mm_interconnect_0|cmd_mux_003|src_payload~19_combout ),
	.src_payload20(\mm_interconnect_0|cmd_mux_003|src_payload~20_combout ),
	.src_payload21(\mm_interconnect_0|cmd_mux_003|src_payload~21_combout ),
	.src_payload22(\mm_interconnect_0|cmd_mux_003|src_payload~22_combout ),
	.src_payload23(\mm_interconnect_0|cmd_mux_003|src_payload~23_combout ),
	.src_payload24(\mm_interconnect_0|cmd_mux_003|src_payload~24_combout ),
	.src_payload25(\mm_interconnect_0|cmd_mux_003|src_payload~25_combout ),
	.src_payload26(\mm_interconnect_0|cmd_mux_003|src_payload~26_combout ),
	.src_payload27(\mm_interconnect_0|cmd_mux_003|src_payload~27_combout ),
	.src_payload28(\mm_interconnect_0|cmd_mux_003|src_payload~28_combout ),
	.src_payload29(\mm_interconnect_0|cmd_mux_003|src_payload~29_combout ),
	.src_payload30(\mm_interconnect_0|cmd_mux_003|src_payload~30_combout ),
	.src_payload31(\mm_interconnect_0|cmd_mux_003|src_payload~31_combout ),
	.clk_clk(\clk_clk~input_o ));

processor_processor_led_pio led_pio(
	.writedata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\cpu|M_st_data[9]~q ,\cpu|M_st_data[8]~q ,\cpu|M_st_data[7]~q ,\cpu|M_st_data[6]~q ,\cpu|M_st_data[5]~q ,\cpu|M_st_data[4]~q ,\cpu|M_st_data[3]~q ,\cpu|M_st_data[2]~q ,\cpu|M_st_data[1]~q ,
\cpu|M_st_data[0]~q }),
	.data_out_0(\led_pio|data_out[0]~q ),
	.data_out_1(\led_pio|data_out[1]~q ),
	.data_out_2(\led_pio|data_out[2]~q ),
	.data_out_3(\led_pio|data_out[3]~q ),
	.data_out_4(\led_pio|data_out[4]~q ),
	.data_out_5(\led_pio|data_out[5]~q ),
	.data_out_6(\led_pio|data_out[6]~q ),
	.data_out_7(\led_pio|data_out[7]~q ),
	.data_out_8(\led_pio|data_out[8]~q ),
	.data_out_9(\led_pio|data_out[9]~q ),
	.reset_n(\rst_controller|r_sync_rst~q ),
	.clr_break_line(\cpu|clr_break_line~q ),
	.d_write(\cpu|d_write~q ),
	.mem_used_1(\mm_interconnect_0|led_pio_s1_agent_rsp_fifo|mem_used[1]~q ),
	.Equal4(\mm_interconnect_0|router|Equal4~0_combout ),
	.wait_latency_counter_1(\mm_interconnect_0|led_pio_s1_translator|wait_latency_counter[1]~q ),
	.wait_latency_counter_0(\mm_interconnect_0|led_pio_s1_translator|wait_latency_counter[0]~q ),
	.M_alu_result_3(\cpu|M_alu_result[3]~q ),
	.M_alu_result_2(\cpu|M_alu_result[2]~q ),
	.readdata_0(\led_pio|readdata[0]~combout ),
	.readdata_8(\led_pio|readdata[8]~combout ),
	.readdata_5(\led_pio|readdata[5]~combout ),
	.readdata_4(\led_pio|readdata[4]~combout ),
	.readdata_6(\led_pio|readdata[6]~combout ),
	.readdata_7(\led_pio|readdata[7]~combout ),
	.readdata_9(\led_pio|readdata[9]~combout ),
	.readdata_3(\led_pio|readdata[3]~combout ),
	.readdata_2(\led_pio|readdata[2]~combout ),
	.readdata_1(\led_pio|readdata[1]~combout ),
	.clk(\clk_clk~input_o ));

processor_processor_mm_interconnect_0 mm_interconnect_0(
	.M_st_data_8(\cpu|M_st_data[8]~q ),
	.M_st_data_9(\cpu|M_st_data[9]~q ),
	.q_a_0(\onchip_mem|the_altsyncram|auto_generated|q_a[0] ),
	.q_a_16(\onchip_mem|the_altsyncram|auto_generated|q_a[16] ),
	.q_a_8(\onchip_mem|the_altsyncram|auto_generated|q_a[8] ),
	.q_a_24(\onchip_mem|the_altsyncram|auto_generated|q_a[24] ),
	.q_a_5(\onchip_mem|the_altsyncram|auto_generated|q_a[5] ),
	.q_a_21(\onchip_mem|the_altsyncram|auto_generated|q_a[21] ),
	.q_a_13(\onchip_mem|the_altsyncram|auto_generated|q_a[13] ),
	.q_a_29(\onchip_mem|the_altsyncram|auto_generated|q_a[29] ),
	.q_a_4(\onchip_mem|the_altsyncram|auto_generated|q_a[4] ),
	.q_a_20(\onchip_mem|the_altsyncram|auto_generated|q_a[20] ),
	.q_a_12(\onchip_mem|the_altsyncram|auto_generated|q_a[12] ),
	.q_a_28(\onchip_mem|the_altsyncram|auto_generated|q_a[28] ),
	.q_a_6(\onchip_mem|the_altsyncram|auto_generated|q_a[6] ),
	.q_a_22(\onchip_mem|the_altsyncram|auto_generated|q_a[22] ),
	.q_a_14(\onchip_mem|the_altsyncram|auto_generated|q_a[14] ),
	.q_a_30(\onchip_mem|the_altsyncram|auto_generated|q_a[30] ),
	.q_a_7(\onchip_mem|the_altsyncram|auto_generated|q_a[7] ),
	.q_a_23(\onchip_mem|the_altsyncram|auto_generated|q_a[23] ),
	.q_a_15(\onchip_mem|the_altsyncram|auto_generated|q_a[15] ),
	.q_a_31(\onchip_mem|the_altsyncram|auto_generated|q_a[31] ),
	.q_a_11(\onchip_mem|the_altsyncram|auto_generated|q_a[11] ),
	.q_a_27(\onchip_mem|the_altsyncram|auto_generated|q_a[27] ),
	.q_a_10(\onchip_mem|the_altsyncram|auto_generated|q_a[10] ),
	.q_a_26(\onchip_mem|the_altsyncram|auto_generated|q_a[26] ),
	.q_a_25(\onchip_mem|the_altsyncram|auto_generated|q_a[25] ),
	.q_a_9(\onchip_mem|the_altsyncram|auto_generated|q_a[9] ),
	.q_a_3(\onchip_mem|the_altsyncram|auto_generated|q_a[3] ),
	.q_a_19(\onchip_mem|the_altsyncram|auto_generated|q_a[19] ),
	.q_a_2(\onchip_mem|the_altsyncram|auto_generated|q_a[2] ),
	.q_a_18(\onchip_mem|the_altsyncram|auto_generated|q_a[18] ),
	.q_a_1(\onchip_mem|the_altsyncram|auto_generated|q_a[1] ),
	.q_a_17(\onchip_mem|the_altsyncram|auto_generated|q_a[17] ),
	.readdata_0(\cpu|the_processor_cpu_nios2_oci|readdata[0]~q ),
	.q_b_0(\jtag_uart|the_processor_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[0] ),
	.Add1(\jtag_uart|Add1~1_sumout ),
	.readdata_16(\cpu|the_processor_cpu_nios2_oci|readdata[16]~q ),
	.M_st_data_16(\cpu|M_st_data[16]~q ),
	.readdata_8(\cpu|the_processor_cpu_nios2_oci|readdata[8]~q ),
	.readdata_24(\cpu|the_processor_cpu_nios2_oci|readdata[24]~q ),
	.readdata_5(\cpu|the_processor_cpu_nios2_oci|readdata[5]~q ),
	.q_b_5(\jtag_uart|the_processor_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[5] ),
	.readdata_21(\cpu|the_processor_cpu_nios2_oci|readdata[21]~q ),
	.M_st_data_21(\cpu|M_st_data[21]~q ),
	.Add11(\jtag_uart|Add1~5_sumout ),
	.readdata_13(\cpu|the_processor_cpu_nios2_oci|readdata[13]~q ),
	.M_st_data_13(\cpu|M_st_data[13]~q ),
	.readdata_29(\cpu|the_processor_cpu_nios2_oci|readdata[29]~q ),
	.readdata_4(\cpu|the_processor_cpu_nios2_oci|readdata[4]~q ),
	.q_b_4(\jtag_uart|the_processor_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[4] ),
	.readdata_20(\cpu|the_processor_cpu_nios2_oci|readdata[20]~q ),
	.M_st_data_20(\cpu|M_st_data[20]~q ),
	.Add12(\jtag_uart|Add1~9_sumout ),
	.readdata_12(\cpu|the_processor_cpu_nios2_oci|readdata[12]~q ),
	.M_st_data_12(\cpu|M_st_data[12]~q ),
	.readdata_28(\cpu|the_processor_cpu_nios2_oci|readdata[28]~q ),
	.readdata_6(\cpu|the_processor_cpu_nios2_oci|readdata[6]~q ),
	.q_b_6(\jtag_uart|the_processor_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[6] ),
	.readdata_22(\cpu|the_processor_cpu_nios2_oci|readdata[22]~q ),
	.M_st_data_22(\cpu|M_st_data[22]~q ),
	.Add13(\jtag_uart|Add1~13_sumout ),
	.readdata_14(\cpu|the_processor_cpu_nios2_oci|readdata[14]~q ),
	.M_st_data_14(\cpu|M_st_data[14]~q ),
	.readdata_30(\cpu|the_processor_cpu_nios2_oci|readdata[30]~q ),
	.readdata_7(\cpu|the_processor_cpu_nios2_oci|readdata[7]~q ),
	.q_b_7(\jtag_uart|the_processor_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[7] ),
	.readdata_23(\cpu|the_processor_cpu_nios2_oci|readdata[23]~q ),
	.M_st_data_23(\cpu|M_st_data[23]~q ),
	.readdata_15(\cpu|the_processor_cpu_nios2_oci|readdata[15]~q ),
	.M_st_data_15(\cpu|M_st_data[15]~q ),
	.readdata_31(\cpu|the_processor_cpu_nios2_oci|readdata[31]~q ),
	.readdata_11(\cpu|the_processor_cpu_nios2_oci|readdata[11]~q ),
	.M_st_data_11(\cpu|M_st_data[11]~q ),
	.readdata_27(\cpu|the_processor_cpu_nios2_oci|readdata[27]~q ),
	.readdata_10(\cpu|the_processor_cpu_nios2_oci|readdata[10]~q ),
	.M_st_data_10(\cpu|M_st_data[10]~q ),
	.readdata_26(\cpu|the_processor_cpu_nios2_oci|readdata[26]~q ),
	.readdata_25(\cpu|the_processor_cpu_nios2_oci|readdata[25]~q ),
	.readdata_9(\cpu|the_processor_cpu_nios2_oci|readdata[9]~q ),
	.q_b_3(\jtag_uart|the_processor_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[3] ),
	.readdata_3(\cpu|the_processor_cpu_nios2_oci|readdata[3]~q ),
	.readdata_19(\cpu|the_processor_cpu_nios2_oci|readdata[19]~q ),
	.M_st_data_19(\cpu|M_st_data[19]~q ),
	.Add14(\jtag_uart|Add1~17_sumout ),
	.q_b_2(\jtag_uart|the_processor_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[2] ),
	.readdata_2(\cpu|the_processor_cpu_nios2_oci|readdata[2]~q ),
	.Add15(\jtag_uart|Add1~21_sumout ),
	.readdata_18(\cpu|the_processor_cpu_nios2_oci|readdata[18]~q ),
	.M_st_data_18(\cpu|M_st_data[18]~q ),
	.q_b_1(\jtag_uart|the_processor_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|FIFOram|q_b[1] ),
	.readdata_1(\cpu|the_processor_cpu_nios2_oci|readdata[1]~q ),
	.readdata_17(\cpu|the_processor_cpu_nios2_oci|readdata[17]~q ),
	.M_st_data_17(\cpu|M_st_data[17]~q ),
	.Add16(\jtag_uart|Add1~25_sumout ),
	.M_st_data_0(\cpu|M_st_data[0]~q ),
	.r_sync_rst(\rst_controller|r_sync_rst~q ),
	.clr_break_line(\cpu|clr_break_line~q ),
	.d_write(\cpu|d_write~q ),
	.mem_used_1(\mm_interconnect_0|led_pio_s1_agent_rsp_fifo|mem_used[1]~q ),
	.M_alu_result_5(\cpu|M_alu_result[5]~q ),
	.M_alu_result_4(\cpu|M_alu_result[4]~q ),
	.M_alu_result_6(\cpu|M_alu_result[6]~q ),
	.M_alu_result_16(\cpu|M_alu_result[16]~q ),
	.M_alu_result_15(\cpu|M_alu_result[15]~q ),
	.M_alu_result_14(\cpu|M_alu_result[14]~q ),
	.M_alu_result_13(\cpu|M_alu_result[13]~q ),
	.Equal1(\mm_interconnect_0|router|Equal1~0_combout ),
	.M_alu_result_12(\cpu|M_alu_result[12]~q ),
	.M_alu_result_11(\cpu|M_alu_result[11]~q ),
	.M_alu_result_10(\cpu|M_alu_result[10]~q ),
	.M_alu_result_9(\cpu|M_alu_result[9]~q ),
	.M_alu_result_8(\cpu|M_alu_result[8]~q ),
	.M_alu_result_7(\cpu|M_alu_result[7]~q ),
	.Equal2(\mm_interconnect_0|router|Equal2~0_combout ),
	.Equal4(\mm_interconnect_0|router|Equal4~0_combout ),
	.wait_latency_counter_1(\mm_interconnect_0|led_pio_s1_translator|wait_latency_counter[1]~q ),
	.wait_latency_counter_0(\mm_interconnect_0|led_pio_s1_translator|wait_latency_counter[0]~q ),
	.M_alu_result_3(\cpu|M_alu_result[3]~q ),
	.M_alu_result_2(\cpu|M_alu_result[2]~q ),
	.M_st_data_1(\cpu|M_st_data[1]~q ),
	.M_st_data_2(\cpu|M_st_data[2]~q ),
	.M_st_data_3(\cpu|M_st_data[3]~q ),
	.M_st_data_4(\cpu|M_st_data[4]~q ),
	.M_st_data_5(\cpu|M_st_data[5]~q ),
	.M_st_data_6(\cpu|M_st_data[6]~q ),
	.M_st_data_7(\cpu|M_st_data[7]~q ),
	.d_read(\cpu|d_read~q ),
	.WideOr1(\mm_interconnect_0|rsp_mux|WideOr1~combout ),
	.read_accepted(\mm_interconnect_0|cpu_data_master_translator|read_accepted~q ),
	.mem_used_11(\mm_interconnect_0|sys_clk_timer_s1_agent_rsp_fifo|mem_used[1]~q ),
	.wait_latency_counter_11(\mm_interconnect_0|sys_clk_timer_s1_translator|wait_latency_counter[1]~q ),
	.wait_latency_counter_01(\mm_interconnect_0|sys_clk_timer_s1_translator|wait_latency_counter[0]~q ),
	.av_waitrequest(\jtag_uart|av_waitrequest~q ),
	.Equal6(\mm_interconnect_0|router|Equal6~0_combout ),
	.saved_grant_0(\mm_interconnect_0|cmd_mux_002|saved_grant[0]~q ),
	.waitrequest(\cpu|the_processor_cpu_nios2_oci|the_processor_cpu_nios2_ocimem|waitrequest~q ),
	.mem_used_12(\mm_interconnect_0|cpu_jtag_debug_module_agent_rsp_fifo|mem_used[1]~q ),
	.saved_grant_01(\mm_interconnect_0|cmd_mux_003|saved_grant[0]~q ),
	.mem_used_13(\mm_interconnect_0|onchip_mem_s1_agent_rsp_fifo|mem_used[1]~q ),
	.read_accepted1(\mm_interconnect_0|cpu_data_master_translator|read_accepted~0_combout ),
	.hbreak_enabled(\cpu|hbreak_enabled~q ),
	.uav_read(\mm_interconnect_0|cpu_data_master_translator|uav_read~0_combout ),
	.src2_valid(\mm_interconnect_0|cmd_demux|src2_valid~2_combout ),
	.saved_grant_1(\mm_interconnect_0|cmd_mux_002|saved_grant[1]~q ),
	.i_read(\cpu|i_read~q ),
	.has_pending_responses(\mm_interconnect_0|cpu_instruction_master_limiter|has_pending_responses~q ),
	.ic_fill_tag_5(\cpu|ic_fill_tag[5]~q ),
	.ic_fill_tag_4(\cpu|ic_fill_tag[4]~q ),
	.ic_fill_tag_3(\cpu|ic_fill_tag[3]~q ),
	.ic_fill_tag_2(\cpu|ic_fill_tag[2]~q ),
	.ic_fill_tag_1(\cpu|ic_fill_tag[1]~q ),
	.ic_fill_tag_0(\cpu|ic_fill_tag[0]~q ),
	.Equal11(\mm_interconnect_0|router_001|Equal1~0_combout ),
	.src0_valid(\mm_interconnect_0|cmd_demux_001|src0_valid~0_combout ),
	.rf_source_valid(\mm_interconnect_0|cpu_jtag_debug_module_agent|rf_source_valid~0_combout ),
	.src3_valid(\mm_interconnect_0|cmd_demux|src3_valid~0_combout ),
	.saved_grant_11(\mm_interconnect_0|cmd_mux_003|saved_grant[1]~q ),
	.last_dest_id_1(\mm_interconnect_0|cpu_instruction_master_limiter|last_dest_id[1]~q ),
	.src1_valid(\mm_interconnect_0|cmd_demux_001|src1_valid~0_combout ),
	.read_latency_shift_reg(\mm_interconnect_0|jtag_uart_avalon_jtag_slave_translator|read_latency_shift_reg~0_combout ),
	.period_l_wr_strobe(\sys_clk_timer|period_l_wr_strobe~0_combout ),
	.src_data_0(\mm_interconnect_0|rsp_mux|src_data[0]~combout ),
	.src_payload(\mm_interconnect_0|rsp_mux|src_payload~1_combout ),
	.src_data_8(\mm_interconnect_0|rsp_mux|src_data[8]~combout ),
	.src_payload1(\mm_interconnect_0|rsp_mux|src_payload~2_combout ),
	.WideOr0(\mm_interconnect_0|cmd_demux_001|WideOr0~0_combout ),
	.nonposted_cmd_accepted(\mm_interconnect_0|cpu_instruction_master_limiter|nonposted_cmd_accepted~combout ),
	.ic_fill_line_5(\cpu|ic_fill_line[5]~q ),
	.src_data_46(\mm_interconnect_0|cmd_mux_002|src_data[46]~combout ),
	.src_data_5(\mm_interconnect_0|rsp_mux|src_data[5]~combout ),
	.src_payload2(\mm_interconnect_0|rsp_mux|src_payload~4_combout ),
	.src_payload3(\mm_interconnect_0|rsp_mux|src_payload~6_combout ),
	.src_payload4(\mm_interconnect_0|rsp_mux|src_payload~7_combout ),
	.src_data_4(\mm_interconnect_0|rsp_mux|src_data[4]~combout ),
	.src_payload5(\mm_interconnect_0|rsp_mux|src_payload~9_combout ),
	.src_payload6(\mm_interconnect_0|rsp_mux|src_payload~11_combout ),
	.src_payload7(\mm_interconnect_0|rsp_mux|src_payload~12_combout ),
	.src_data_6(\mm_interconnect_0|rsp_mux|src_data[6]~combout ),
	.src_payload8(\mm_interconnect_0|rsp_mux|src_payload~14_combout ),
	.src_payload9(\mm_interconnect_0|rsp_mux|src_payload~16_combout ),
	.src_payload10(\mm_interconnect_0|rsp_mux|src_payload~17_combout ),
	.src_data_7(\mm_interconnect_0|rsp_mux|src_data[7]~combout ),
	.src_payload11(\mm_interconnect_0|rsp_mux|src_payload~18_combout ),
	.src_payload12(\mm_interconnect_0|rsp_mux|src_payload~20_combout ),
	.src_payload13(\mm_interconnect_0|rsp_mux|src_payload~21_combout ),
	.ien_AE(\jtag_uart|ien_AE~q ),
	.av_readdata_9(\jtag_uart|av_readdata[9]~combout ),
	.ien_AF(\jtag_uart|ien_AF~q ),
	.av_readdata_8(\jtag_uart|av_readdata[8]~0_combout ),
	.src_payload14(\mm_interconnect_0|rsp_mux|src_payload~22_combout ),
	.src_payload15(\mm_interconnect_0|rsp_mux|src_payload~23_combout ),
	.src_payload16(\mm_interconnect_0|rsp_mux|src_payload~25_combout ),
	.src_payload17(\mm_interconnect_0|rsp_mux|src_payload~26_combout ),
	.src_payload18(\mm_interconnect_0|rsp_mux|src_payload~27_combout ),
	.src_data_9(\mm_interconnect_0|rsp_mux|src_data[9]~combout ),
	.src_data_3(\mm_interconnect_0|rsp_mux|src_data[3]~combout ),
	.src_payload19(\mm_interconnect_0|rsp_mux|src_payload~29_combout ),
	.src_data_2(\mm_interconnect_0|rsp_mux|src_data[2]~combout ),
	.src_payload20(\mm_interconnect_0|rsp_mux|src_payload~30_combout ),
	.src_data_1(\mm_interconnect_0|rsp_mux|src_data[1]~combout ),
	.src_payload21(\mm_interconnect_0|rsp_mux|src_payload~32_combout ),
	.b_full(\jtag_uart|the_processor_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|b_full~q ),
	.ic_fill_line_0(\cpu|ic_fill_line[0]~q ),
	.ic_fill_line_1(\cpu|ic_fill_line[1]~q ),
	.ic_fill_line_2(\cpu|ic_fill_line[2]~q ),
	.ic_fill_line_3(\cpu|ic_fill_line[3]~q ),
	.ic_fill_line_4(\cpu|ic_fill_line[4]~q ),
	.src_payload22(\mm_interconnect_0|cmd_mux_003|src_payload~0_combout ),
	.ic_fill_ap_offset_0(\cpu|ic_fill_ap_offset[0]~q ),
	.src_data_38(\mm_interconnect_0|cmd_mux_003|src_data[38]~combout ),
	.ic_fill_ap_offset_1(\cpu|ic_fill_ap_offset[1]~q ),
	.src_data_39(\mm_interconnect_0|cmd_mux_003|src_data[39]~combout ),
	.ic_fill_ap_offset_2(\cpu|ic_fill_ap_offset[2]~q ),
	.src_data_40(\mm_interconnect_0|cmd_mux_003|src_data[40]~combout ),
	.src_data_41(\mm_interconnect_0|cmd_mux_003|src_data[41]~combout ),
	.src_data_42(\mm_interconnect_0|cmd_mux_003|src_data[42]~combout ),
	.src_data_43(\mm_interconnect_0|cmd_mux_003|src_data[43]~combout ),
	.src_data_44(\mm_interconnect_0|cmd_mux_003|src_data[44]~combout ),
	.src_data_45(\mm_interconnect_0|cmd_mux_003|src_data[45]~combout ),
	.src_data_461(\mm_interconnect_0|cmd_mux_003|src_data[46]~combout ),
	.src_data_47(\mm_interconnect_0|cmd_mux_003|src_data[47]~combout ),
	.src_data_48(\mm_interconnect_0|cmd_mux_003|src_data[48]~combout ),
	.src_data_49(\mm_interconnect_0|cmd_mux_003|src_data[49]~combout ),
	.src_data_50(\mm_interconnect_0|cmd_mux_003|src_data[50]~combout ),
	.M_mem_byte_en_0(\cpu|M_mem_byte_en[0]~q ),
	.src_data_32(\mm_interconnect_0|cmd_mux_003|src_data[32]~combout ),
	.readdata_01(\switches_pio|readdata[0]~q ),
	.readdata_02(\led_pio|readdata[0]~combout ),
	.read_0(\jtag_uart|read_0~q ),
	.readdata_03(\sys_clk_timer|readdata[0]~q ),
	.counter_reg_bit_0(\jtag_uart|the_processor_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[0]~q ),
	.src_payload23(\mm_interconnect_0|cmd_mux_003|src_payload~1_combout ),
	.M_mem_byte_en_2(\cpu|M_mem_byte_en[2]~q ),
	.src_data_34(\mm_interconnect_0|cmd_mux_003|src_data[34]~combout ),
	.src_payload24(\mm_interconnect_0|cmd_mux_003|src_payload~2_combout ),
	.M_mem_byte_en_1(\cpu|M_mem_byte_en[1]~q ),
	.src_data_33(\mm_interconnect_0|cmd_mux_003|src_data[33]~combout ),
	.readdata_81(\led_pio|readdata[8]~combout ),
	.readdata_82(\sys_clk_timer|readdata[8]~q ),
	.readdata_83(\switches_pio|readdata[8]~q ),
	.M_st_data_24(\cpu|M_st_data[24]~q ),
	.src_payload25(\mm_interconnect_0|cmd_mux_003|src_payload~3_combout ),
	.M_mem_byte_en_3(\cpu|M_mem_byte_en[3]~q ),
	.src_data_35(\mm_interconnect_0|cmd_mux_003|src_data[35]~combout ),
	.src_payload26(\mm_interconnect_0|cmd_mux_002|src_payload~0_combout ),
	.src_data_381(\mm_interconnect_0|cmd_mux_002|src_data[38]~combout ),
	.src_data_411(\mm_interconnect_0|cmd_mux_002|src_data[41]~combout ),
	.src_data_401(\mm_interconnect_0|cmd_mux_002|src_data[40]~combout ),
	.src_data_391(\mm_interconnect_0|cmd_mux_002|src_data[39]~combout ),
	.src_data_451(\mm_interconnect_0|cmd_mux_002|src_data[45]~combout ),
	.src_data_441(\mm_interconnect_0|cmd_mux_002|src_data[44]~combout ),
	.src_data_431(\mm_interconnect_0|cmd_mux_002|src_data[43]~combout ),
	.src_data_421(\mm_interconnect_0|cmd_mux_002|src_data[42]~combout ),
	.src_payload27(\mm_interconnect_0|cmd_mux_002|src_payload~1_combout ),
	.src_payload28(\mm_interconnect_0|cmd_mux_003|src_payload~4_combout ),
	.readdata_51(\switches_pio|readdata[5]~q ),
	.readdata_52(\led_pio|readdata[5]~combout ),
	.readdata_53(\sys_clk_timer|readdata[5]~q ),
	.src_payload29(\mm_interconnect_0|cmd_mux_003|src_payload~5_combout ),
	.counter_reg_bit_5(\jtag_uart|the_processor_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[5]~q ),
	.src_payload30(\mm_interconnect_0|cmd_mux_003|src_payload~6_combout ),
	.b_full1(\jtag_uart|the_processor_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|b_full~q ),
	.readdata_131(\sys_clk_timer|readdata[13]~q ),
	.M_st_data_29(\cpu|M_st_data[29]~q ),
	.src_payload31(\mm_interconnect_0|cmd_mux_003|src_payload~7_combout ),
	.src_payload32(\mm_interconnect_0|cmd_mux_003|src_payload~8_combout ),
	.readdata_41(\switches_pio|readdata[4]~q ),
	.readdata_42(\led_pio|readdata[4]~combout ),
	.readdata_43(\sys_clk_timer|readdata[4]~q ),
	.src_payload33(\mm_interconnect_0|cmd_mux_003|src_payload~9_combout ),
	.counter_reg_bit_4(\jtag_uart|the_processor_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[4]~q ),
	.src_payload34(\mm_interconnect_0|cmd_mux_003|src_payload~10_combout ),
	.b_non_empty(\jtag_uart|the_processor_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|b_non_empty~q ),
	.readdata_121(\sys_clk_timer|readdata[12]~q ),
	.M_st_data_28(\cpu|M_st_data[28]~q ),
	.src_payload35(\mm_interconnect_0|cmd_mux_003|src_payload~11_combout ),
	.src_payload36(\mm_interconnect_0|cmd_mux_003|src_payload~12_combout ),
	.readdata_61(\switches_pio|readdata[6]~q ),
	.readdata_62(\led_pio|readdata[6]~combout ),
	.readdata_63(\sys_clk_timer|readdata[6]~q ),
	.src_payload37(\mm_interconnect_0|cmd_mux_003|src_payload~13_combout ),
	.src_payload38(\mm_interconnect_0|cmd_mux_003|src_payload~14_combout ),
	.woverflow(\jtag_uart|woverflow~q ),
	.readdata_141(\sys_clk_timer|readdata[14]~q ),
	.M_st_data_30(\cpu|M_st_data[30]~q ),
	.src_payload39(\mm_interconnect_0|cmd_mux_003|src_payload~15_combout ),
	.src_payload40(\mm_interconnect_0|cmd_mux_003|src_payload~16_combout ),
	.readdata_71(\switches_pio|readdata[7]~q ),
	.readdata_72(\led_pio|readdata[7]~combout ),
	.readdata_73(\sys_clk_timer|readdata[7]~q ),
	.src_payload41(\mm_interconnect_0|cmd_mux_003|src_payload~17_combout ),
	.src_payload42(\mm_interconnect_0|cmd_mux_003|src_payload~18_combout ),
	.rvalid(\jtag_uart|rvalid~q ),
	.readdata_151(\sys_clk_timer|readdata[15]~q ),
	.M_st_data_31(\cpu|M_st_data[31]~q ),
	.src_payload43(\mm_interconnect_0|cmd_mux_003|src_payload~19_combout ),
	.src_payload44(\mm_interconnect_0|cmd_mux_003|src_payload~20_combout ),
	.readdata_111(\sys_clk_timer|readdata[11]~q ),
	.M_st_data_27(\cpu|M_st_data[27]~q ),
	.src_payload45(\mm_interconnect_0|cmd_mux_003|src_payload~21_combout ),
	.src_payload46(\mm_interconnect_0|cmd_mux_003|src_payload~22_combout ),
	.ac(\jtag_uart|ac~q ),
	.readdata_101(\sys_clk_timer|readdata[10]~q ),
	.M_st_data_26(\cpu|M_st_data[26]~q ),
	.src_payload47(\mm_interconnect_0|cmd_mux_003|src_payload~23_combout ),
	.M_st_data_25(\cpu|M_st_data[25]~q ),
	.src_payload48(\mm_interconnect_0|cmd_mux_003|src_payload~24_combout ),
	.src_payload49(\mm_interconnect_0|cmd_mux_003|src_payload~25_combout ),
	.readdata_91(\led_pio|readdata[9]~combout ),
	.readdata_92(\sys_clk_timer|readdata[9]~q ),
	.readdata_93(\switches_pio|readdata[9]~q ),
	.src_payload50(\mm_interconnect_0|cmd_mux_003|src_payload~26_combout ),
	.readdata_32(\led_pio|readdata[3]~combout ),
	.readdata_33(\sys_clk_timer|readdata[3]~q ),
	.readdata_34(\switches_pio|readdata[3]~q ),
	.src_payload51(\mm_interconnect_0|cmd_mux_003|src_payload~27_combout ),
	.counter_reg_bit_3(\jtag_uart|the_processor_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[3]~q ),
	.src_payload52(\mm_interconnect_0|cmd_mux_003|src_payload~28_combout ),
	.readdata_210(\led_pio|readdata[2]~combout ),
	.readdata_211(\sys_clk_timer|readdata[2]~q ),
	.readdata_212(\switches_pio|readdata[2]~q ),
	.counter_reg_bit_2(\jtag_uart|the_processor_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[2]~q ),
	.src_payload53(\mm_interconnect_0|cmd_mux_003|src_payload~29_combout ),
	.src_payload54(\mm_interconnect_0|cmd_mux_003|src_payload~30_combout ),
	.readdata_110(\led_pio|readdata[1]~combout ),
	.readdata_112(\sys_clk_timer|readdata[1]~q ),
	.readdata_113(\switches_pio|readdata[1]~q ),
	.src_payload55(\mm_interconnect_0|cmd_mux_003|src_payload~31_combout ),
	.counter_reg_bit_1(\jtag_uart|the_processor_jtag_uart_scfifo_r|rfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[1]~q ),
	.src_payload56(\mm_interconnect_0|cmd_mux_002|src_payload~2_combout ),
	.src_data_321(\mm_interconnect_0|cmd_mux_002|src_data[32]~combout ),
	.WideOr11(\mm_interconnect_0|rsp_mux_001|WideOr1~combout ),
	.src_data_24(\mm_interconnect_0|rsp_mux_001|src_data[24]~combout ),
	.src_data_01(\mm_interconnect_0|rsp_mux_001|src_data[0]~combout ),
	.src_data_11(\mm_interconnect_0|rsp_mux_001|src_data[1]~combout ),
	.src_data_21(\mm_interconnect_0|rsp_mux_001|src_data[2]~combout ),
	.src_data_31(\mm_interconnect_0|rsp_mux_001|src_data[3]~combout ),
	.src_data_410(\mm_interconnect_0|rsp_mux_001|src_data[4]~combout ),
	.src_data_51(\mm_interconnect_0|rsp_mux_001|src_data[5]~combout ),
	.src_data_22(\mm_interconnect_0|rsp_mux_001|src_data[22]~combout ),
	.src_data_23(\mm_interconnect_0|rsp_mux_001|src_data[23]~combout ),
	.src_data_25(\mm_interconnect_0|rsp_mux_001|src_data[25]~combout ),
	.src_data_26(\mm_interconnect_0|rsp_mux_001|src_data[26]~combout ),
	.src_data_14(\mm_interconnect_0|rsp_mux_001|src_data[14]~combout ),
	.src_data_12(\mm_interconnect_0|rsp_mux_001|src_data[12]~combout ),
	.src_data_111(\mm_interconnect_0|rsp_mux_001|src_data[11]~combout ),
	.src_data_16(\mm_interconnect_0|rsp_mux_001|src_data[16]~combout ),
	.src_data_15(\mm_interconnect_0|rsp_mux_001|src_data[15]~combout ),
	.src_data_13(\mm_interconnect_0|rsp_mux_001|src_data[13]~combout ),
	.src_data_211(\mm_interconnect_0|rsp_mux_001|src_data[21]~combout ),
	.src_data_29(\mm_interconnect_0|rsp_mux_001|src_data[29]~combout ),
	.src_data_27(\mm_interconnect_0|rsp_mux_001|src_data[27]~combout ),
	.src_data_28(\mm_interconnect_0|rsp_mux_001|src_data[28]~combout ),
	.src_data_30(\mm_interconnect_0|rsp_mux_001|src_data[30]~combout ),
	.src_data_311(\mm_interconnect_0|rsp_mux_001|src_data[31]~combout ),
	.src_data_10(\mm_interconnect_0|rsp_mux_001|src_data[10]~combout ),
	.src_data_61(\mm_interconnect_0|rsp_mux_001|src_data[6]~combout ),
	.src_data_81(\mm_interconnect_0|rsp_mux_001|src_data[8]~combout ),
	.src_payload57(\mm_interconnect_0|cmd_mux_002|src_payload~3_combout ),
	.src_data_71(\mm_interconnect_0|rsp_mux_001|src_data[7]~combout ),
	.src_data_20(\mm_interconnect_0|rsp_mux_001|src_data[20]~combout ),
	.src_data_19(\mm_interconnect_0|rsp_mux_001|src_data[19]~combout ),
	.src_data_18(\mm_interconnect_0|rsp_mux_001|src_data[18]~combout ),
	.src_data_17(\mm_interconnect_0|rsp_mux_001|src_data[17]~combout ),
	.src_data_91(\mm_interconnect_0|rsp_mux_001|src_data[9]~combout ),
	.src_payload58(\mm_interconnect_0|cmd_mux_002|src_payload~4_combout ),
	.src_payload59(\mm_interconnect_0|cmd_mux_002|src_payload~5_combout ),
	.src_data_341(\mm_interconnect_0|cmd_mux_002|src_data[34]~combout ),
	.src_payload60(\mm_interconnect_0|cmd_mux_002|src_payload~6_combout ),
	.src_data_331(\mm_interconnect_0|cmd_mux_002|src_data[33]~combout ),
	.src_payload61(\mm_interconnect_0|cmd_mux_002|src_payload~7_combout ),
	.src_data_351(\mm_interconnect_0|cmd_mux_002|src_data[35]~combout ),
	.src_payload62(\mm_interconnect_0|cmd_mux_002|src_payload~8_combout ),
	.src_payload63(\mm_interconnect_0|cmd_mux_002|src_payload~9_combout ),
	.src_payload64(\mm_interconnect_0|cmd_mux_002|src_payload~10_combout ),
	.src_payload65(\mm_interconnect_0|cmd_mux_002|src_payload~11_combout ),
	.src_payload66(\mm_interconnect_0|cmd_mux_002|src_payload~12_combout ),
	.src_payload67(\mm_interconnect_0|cmd_mux_002|src_payload~13_combout ),
	.src_payload68(\mm_interconnect_0|cmd_mux_002|src_payload~14_combout ),
	.src_payload69(\mm_interconnect_0|cmd_mux_002|src_payload~15_combout ),
	.src_payload70(\mm_interconnect_0|cmd_mux_002|src_payload~16_combout ),
	.src_payload71(\mm_interconnect_0|cmd_mux_002|src_payload~17_combout ),
	.src_payload72(\mm_interconnect_0|cmd_mux_002|src_payload~18_combout ),
	.src_payload73(\mm_interconnect_0|cmd_mux_002|src_payload~19_combout ),
	.src_payload74(\mm_interconnect_0|cmd_mux_002|src_payload~20_combout ),
	.src_payload75(\mm_interconnect_0|cmd_mux_002|src_payload~21_combout ),
	.src_payload76(\mm_interconnect_0|cmd_mux_002|src_payload~22_combout ),
	.src_payload77(\mm_interconnect_0|cmd_mux_002|src_payload~23_combout ),
	.src_payload78(\mm_interconnect_0|cmd_mux_002|src_payload~24_combout ),
	.src_payload79(\mm_interconnect_0|cmd_mux_002|src_payload~25_combout ),
	.src_payload80(\mm_interconnect_0|cmd_mux_002|src_payload~26_combout ),
	.src_payload81(\mm_interconnect_0|cmd_mux_002|src_payload~27_combout ),
	.src_payload82(\mm_interconnect_0|cmd_mux_002|src_payload~28_combout ),
	.src_payload83(\mm_interconnect_0|cmd_mux_002|src_payload~29_combout ),
	.src_payload84(\mm_interconnect_0|cmd_mux_002|src_payload~30_combout ),
	.src_payload85(\mm_interconnect_0|cmd_mux_002|src_payload~31_combout ),
	.src_payload86(\mm_interconnect_0|cmd_mux_002|src_payload~32_combout ),
	.GND_port(\~GND~combout ),
	.clk_clk(\clk_clk~input_o ));

processor_altera_reset_controller rst_controller(
	.r_sync_rst1(\rst_controller|r_sync_rst~q ),
	.r_early_rst1(\rst_controller|r_early_rst~q ),
	.altera_reset_synchronizer_int_chain_1(\rst_controller|alt_rst_req_sync_uq1|altera_reset_synchronizer_int_chain[1]~0_combout ),
	.clk_clk(\clk_clk~input_o ),
	.reset_reset_n(\reset_reset_n~input_o ));

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~1_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_1[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~3_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_1[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_1[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_1[3] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~3_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~5_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~6_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~5_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][1] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0 .lut_mask = 64'hFEFEFEFEFEFEFEFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~1 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\altera_internal_jtag~TDIUTAP ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~1 .lut_mask = 64'hEDDEFFFFFFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~1 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2 .lut_mask = 64'h7FBFFFFFFFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~3 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\altera_internal_jtag~TDIUTAP ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~3 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~3 .lut_mask = 64'hFFFFB77BFFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~3 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~5_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~6_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~3 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~3 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~3 .lut_mask = 64'h4747474747474747;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~3 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~14 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~14 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~14 .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~14 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~4 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~4 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~4 .lut_mask = 64'hFFFFEFFFFFFFFFEF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~4 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~5 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~14_combout ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~4_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~5 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~5 .lut_mask = 64'hFFF7FFFFFFF7FFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~5 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~7_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~6_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][1] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~6 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~6 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~6 .lut_mask = 64'h4747474747474747;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~6 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~5 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~5 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~5 .lut_mask = 64'h2727272727272727;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~5 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~6 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~14_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~6 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~6 .lut_mask = 64'hFFFFFFFF7FFFF7FF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~6 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~7 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][1]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~7 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~7 .lut_mask = 64'h2727272727272727;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~7 .shared_arith = "off";

assign \clk_clk~input_o  = clk_clk;

assign \switches_pio_external_connection_export[0]~input_o  = switches_pio_external_connection_export[0];

assign \switches_pio_external_connection_export[8]~input_o  = switches_pio_external_connection_export[8];

assign \switches_pio_external_connection_export[5]~input_o  = switches_pio_external_connection_export[5];

assign \switches_pio_external_connection_export[4]~input_o  = switches_pio_external_connection_export[4];

assign \switches_pio_external_connection_export[6]~input_o  = switches_pio_external_connection_export[6];

assign \switches_pio_external_connection_export[7]~input_o  = switches_pio_external_connection_export[7];

assign \switches_pio_external_connection_export[9]~input_o  = switches_pio_external_connection_export[9];

assign \switches_pio_external_connection_export[3]~input_o  = switches_pio_external_connection_export[3];

assign \switches_pio_external_connection_export[2]~input_o  = switches_pio_external_connection_export[2];

assign \switches_pio_external_connection_export[1]~input_o  = switches_pio_external_connection_export[1];

assign \reset_reset_n~input_o  = reset_reset_n;

assign led_pio_external_connection_export[0] = \led_pio|data_out[0]~q ;

assign led_pio_external_connection_export[1] = \led_pio|data_out[1]~q ;

assign led_pio_external_connection_export[2] = \led_pio|data_out[2]~q ;

assign led_pio_external_connection_export[3] = \led_pio|data_out[3]~q ;

assign led_pio_external_connection_export[4] = \led_pio|data_out[4]~q ;

assign led_pio_external_connection_export[5] = \led_pio|data_out[5]~q ;

assign led_pio_external_connection_export[6] = \led_pio|data_out[6]~q ;

assign led_pio_external_connection_export[7] = \led_pio|data_out[7]~q ;

assign led_pio_external_connection_export[8] = \led_pio|data_out[8]~q ;

assign led_pio_external_connection_export[9] = \led_pio|data_out[9]~q ;

assign altera_reserved_tdo = \altera_internal_jtag~TDO ;

assign \altera_reserved_tms~input_o  = altera_reserved_tms;

assign \altera_reserved_tck~input_o  = altera_reserved_tck;

assign \altera_reserved_tdi~input_o  = altera_reserved_tdi;

cyclonev_jtag altera_internal_jtag(
	.tms(\altera_reserved_tms~input_o ),
	.tck(\altera_reserved_tck~input_o ),
	.tdi(\altera_reserved_tdi~input_o ),
	.tdoutap(gnd),
	.tdouser(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~q ),
	.tdo(\altera_internal_jtag~TDO ),
	.tmsutap(\altera_internal_jtag~TMSUTAP ),
	.tckutap(\altera_internal_jtag~TCKUTAP ),
	.tdiutap(\altera_internal_jtag~TDIUTAP ),
	.shiftuser(),
	.clkdruser(),
	.updateuser(),
	.runidleuser(),
	.usr1user());

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0 .lut_mask = 64'h7777777777777777;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~1 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~1 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~1 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~2 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~2 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~2 .lut_mask = 64'h6666666666666666;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~2 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~0 .lut_mask = 64'h9696969696969696;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~0 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~0 .lut_mask = 64'hFFFBFFFBFFFBFFFB;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~6 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~6 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~6 .lut_mask = 64'h7777777777777777;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~6 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~7 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~7 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~7 .lut_mask = 64'h7777777777777777;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~7 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~4 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~4 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~4 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~4 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~5 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~5 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~5 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~5 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~9 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~9 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~9 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~9 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~12 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~12 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~12 .lut_mask = 64'h7777777777777777;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~12 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~13 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~13 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~13 .lut_mask = 64'h7777777777777777;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~13 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~10 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~10 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~10 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~10 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~11 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~11 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~11 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~11 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~1 .lut_mask = 64'hBFFFBFFFBFFFBFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~1 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~2 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~2 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~2 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~2 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~3 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~3 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~3 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~3 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0 .lut_mask = 64'h7777777777777777;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\altera_internal_jtag~TDIUTAP ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~0_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~1 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~1 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~1_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0 .lut_mask = 64'hFFFFFFFEFFFFFFFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal1~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal1~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal1~0 .lut_mask = 64'hFFFFFFEFFFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal1~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal1~0_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg .power_up = "low";

cyclonev_lcell_comb \~GND (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\~GND~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \~GND .extended_lut = "off";
defparam \~GND .lut_mask = 64'h0000000000000000;
defparam \~GND .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~8 (
	.dataa(!\rst_controller|alt_rst_req_sync_uq1|altera_reset_synchronizer_int_chain[1]~0_combout ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datac(!\~GND~combout ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.dataf(!\altera_internal_jtag~TDIUTAP ),
	.datag(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~8 .extended_lut = "on";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~8 .lut_mask = 64'hEFFEFAFCEFFEFAFC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~8 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~5 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~5 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~5 .lut_mask = 64'h96FFFFFF96FFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~5 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~5_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~6 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~6 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~6 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~6 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~4 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.datad(!\cpu|the_processor_cpu_nios2_oci|the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_tck|ir_out[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~4 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~4 .lut_mask = 64'h47FF47FF47FF47FF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~4 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~4_combout ),
	.asdata(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~2_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg~3 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg~3 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg~3 .lut_mask = 64'hFFFFFFDFFFFFFFDF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg~3 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg~3_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~1 .lut_mask = 64'hFFFFFFACFFFFFFAC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~1 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~2 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~2 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~2 .lut_mask = 64'hDF1FDF1FDF1FDF1F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~2 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~6_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~2_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~7 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~7 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~7 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~7 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~7_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~2_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~3 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~3 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~3 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~3 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~3_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~2_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal11~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal11~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal11~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal11~0 .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal11~0 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal11~0_combout ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~0 .lut_mask = 64'hFDDFFFFFDFFDFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~0_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~1 .lut_mask = 64'hFFF7FFF7FFF7FFF7;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~1 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~2 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~2 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~2 .lut_mask = 64'hCF5FFFFFCF5FFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~2 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~2_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg_proc~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg_proc~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg_proc~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg_proc~0 .lut_mask = 64'h7777777777777777;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg_proc~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg_proc~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~8_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~1 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~1 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~2 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~2 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~2 .lut_mask = 64'hEFFFEFFFEFFFEFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~2 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~3 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~3 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~3 .lut_mask = 64'h2727272727272727;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~3 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~4 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8_combout ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~1_combout ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~2_combout ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~3_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~4 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~4 .lut_mask = 64'h6F9F9F6FFFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~4 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~4_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0 .lut_mask = 64'hEFDFDFEFFFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~0 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~0 .lut_mask = 64'hF7FFFFFFF7FFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~0 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~1 .lut_mask = 64'hF7FFFFF7FFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~1 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~2 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0_combout ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~0_combout ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~2 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~2 .lut_mask = 64'h7FFFF7FFFFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~2 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~2_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datab(!\cpu|the_processor_cpu_nios2_oci|the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_tck|ir_out[0]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~0 .lut_mask = 64'hB77BFFFFB77BFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~0_combout ),
	.asdata(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~2_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_tdo_sel_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_tdo_sel_reg[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_tdo_sel_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_tdo_sel_reg[1] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_tdo_sel_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_tdo_sel_reg[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_tdo_sel_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_tdo_sel_reg[0] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datac(!\jtag_uart|processor_jtag_uart_alt_jtag_atlantic|tdo~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_tdo_sel_reg[1]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_tdo_sel_reg[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~0 .lut_mask = 64'hFF3F7F7FFF3F7F7F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~0 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal .lut_mask = 64'h7777777777777777;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~5 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~5 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~5 .lut_mask = 64'hFFAAAAFFAAFFFFAA;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~5 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1 .lut_mask = 64'hFFFFFFDFFFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~1 .lut_mask = 64'hF7FFFFFFF7FFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~1 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~2 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~2 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~2 .lut_mask = 64'hEBBEBEEBBEEBEBBE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~2 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~0 .lut_mask = 64'hFBFEFEFBFEFBFBFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~4 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~4 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~4 .lut_mask = 64'hFFFFFEFFFFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~4 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~3 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~3 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~3 .lut_mask = 64'hAAFFFFAAAAFFFFAA;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~3 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~5 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~5 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~5 .lut_mask = 64'hFFFFFEFFFFFFFEFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~5 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~8 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ),
	.datac(!\altera_internal_jtag~TDIUTAP ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datag(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~8 .extended_lut = "on";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~8 .lut_mask = 64'hFFF7FFF7FFF7FFF7;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~8 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~2 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~2 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~2 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~2 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~2_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[3] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~6 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~6 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~6 .lut_mask = 64'hDF8FDF8FDF8FDF8F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~6 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~7 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~5_combout ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[3]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~6_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~7 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~7 .lut_mask = 64'hD8FFFFFFFFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~7 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~2_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~3 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~3 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~3 .lut_mask = 64'h7777777777777777;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~3 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~4 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~3_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~4 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~4 .lut_mask = 64'hFFFFFFFFDF8FFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~4 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~2_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~0 .lut_mask = 64'h6996699669966996;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~0 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~1 .lut_mask = 64'hF7B3FFFFF7B3FFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~1 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~2_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal11~0_combout ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~1 .lut_mask = 64'hFFFEFFFFFFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~1 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~2 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.datad(!\jtag_uart|processor_jtag_uart_alt_jtag_atlantic|tdo~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_tdo_sel_reg[1]~q ),
	.dataf(!\cpu|the_processor_cpu_nios2_oci|the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_tck|sr[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~2 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~2 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~2 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~0 (
	.dataa(!\altera_internal_jtag~TDIUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~0 .lut_mask = 64'h4747474747474747;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~3 (
	.dataa(!\altera_internal_jtag~TDIUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~3 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~3 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~3 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[3] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~2 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~2 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~2 .lut_mask = 64'h7777777777777777;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~2 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[2] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~1 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~1 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[1] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~0 .lut_mask = 64'h7777777777777777;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[0] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0 .lut_mask = 64'h7777777777777777;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~4 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datae(gnd),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~4 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~4 .lut_mask = 64'hFF00FF00FFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~4 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~1 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~1 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~3 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datae(gnd),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~3 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~3 .lut_mask = 64'h0FF00FF0FFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~3 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.datab(gnd),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datae(gnd),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~0 .lut_mask = 64'hA55AA55AFFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~5 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.datab(gnd),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~5 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~5 .lut_mask = 64'h5AA5A55AFFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~5 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~2 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~2 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~2 .lut_mask = 64'h96696996FFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~2 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~0 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~0 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~1 .lut_mask = 64'hFEEFEFFEFEEFEFFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~1 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~4 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~4 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~4 .lut_mask = 64'hBEEBEBBEBEEBEBBE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~4 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~6 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~6 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~6 .lut_mask = 64'h9669699696696996;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~6 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~8 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~8 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~8 .lut_mask = 64'h9669699696696996;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~8 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal11~0_combout ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0 .lut_mask = 64'hDFFFFFFFFFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\altera_internal_jtag~TDIUTAP ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0 .lut_mask = 64'hFBFFFFFFFBFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[3] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~9 (
	.dataa(!\altera_internal_jtag~TDIUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0_combout ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~0_combout ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~8_combout ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[3]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~9 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~9 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~9 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~3 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~3 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~3 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~3 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~3_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[2] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~7 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0_combout ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~0_combout ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~6_combout ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[2]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~7 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~7 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~7 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~3_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[1] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~5 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0_combout ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~0_combout ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~4_combout ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~5 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~5 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~5 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~3_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~2 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0_combout ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~0_combout ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~1_combout ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~2 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~2 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~2 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~3_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~3 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~3 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~3 .lut_mask = 64'h4747474747474747;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~3 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~4 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~4 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~4 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~4 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~5 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~5 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~5 .lut_mask = 64'hFFFFFFFFFFFFBFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~5 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~6 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~3_combout ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~4_combout ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~5_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~6 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~6 .lut_mask = 64'hFFFFFFFFFFFBFFFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~6 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~7 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~0_combout ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~1_combout ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~2_combout ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~6_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~7 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~7 .lut_mask = 64'hFFFF7FFFFFFF7FFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~7 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo (
	.clk(!\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo .power_up = "low";

cyclonev_lcell_comb \auto_hub|~GND (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|~GND~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|~GND .extended_lut = "off";
defparam \auto_hub|~GND .lut_mask = 64'h0000000000000000;
defparam \auto_hub|~GND .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~_wirecell (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~_wirecell_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~_wirecell .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~_wirecell .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~_wirecell (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~_wirecell_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~_wirecell .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~_wirecell .shared_arith = "off";

endmodule

module processor_altera_reset_controller (
	r_sync_rst1,
	r_early_rst1,
	altera_reset_synchronizer_int_chain_1,
	clk_clk,
	reset_reset_n)/* synthesis synthesis_greybox=1 */;
output 	r_sync_rst1;
output 	r_early_rst1;
output 	altera_reset_synchronizer_int_chain_1;
input 	clk_clk;
input 	reset_reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \alt_rst_req_sync_uq1|altera_reset_synchronizer_int_chain_out~q ;
wire \alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ;
wire \altera_reset_synchronizer_int_chain[0]~q ;
wire \altera_reset_synchronizer_int_chain[1]~q ;
wire \altera_reset_synchronizer_int_chain[2]~q ;
wire \altera_reset_synchronizer_int_chain[3]~q ;
wire \altera_reset_synchronizer_int_chain[4]~0_combout ;
wire \altera_reset_synchronizer_int_chain[4]~q ;
wire \r_sync_rst_chain[3]~q ;
wire \r_sync_rst_chain~1_combout ;
wire \r_sync_rst_chain[2]~q ;
wire \r_sync_rst_chain~0_combout ;
wire \r_sync_rst_chain[1]~q ;
wire \WideOr0~0_combout ;
wire \always2~0_combout ;


processor_altera_reset_synchronizer alt_rst_req_sync_uq1(
	.altera_reset_synchronizer_int_chain_out1(\alt_rst_req_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.altera_reset_synchronizer_int_chain_1(altera_reset_synchronizer_int_chain_1),
	.clk(clk_clk));

processor_altera_reset_synchronizer_1 alt_rst_sync_uq1(
	.altera_reset_synchronizer_int_chain_out1(\alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.clk(clk_clk),
	.reset_reset_n(reset_reset_n));

dffeas r_sync_rst(
	.clk(clk_clk),
	.d(\WideOr0~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(r_sync_rst1),
	.prn(vcc));
defparam r_sync_rst.is_wysiwyg = "true";
defparam r_sync_rst.power_up = "low";

dffeas r_early_rst(
	.clk(clk_clk),
	.d(\always2~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(r_early_rst1),
	.prn(vcc));
defparam r_early_rst.is_wysiwyg = "true";
defparam r_early_rst.power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[0] (
	.clk(clk_clk),
	.d(\alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[0]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[0] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[0] .power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[1] (
	.clk(clk_clk),
	.d(\altera_reset_synchronizer_int_chain[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[1]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[1] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[1] .power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[2] (
	.clk(clk_clk),
	.d(\altera_reset_synchronizer_int_chain[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[2]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[2] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[2] .power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[3] (
	.clk(clk_clk),
	.d(\altera_reset_synchronizer_int_chain[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[3]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[3] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[3] .power_up = "low";

cyclonev_lcell_comb \altera_reset_synchronizer_int_chain[4]~0 (
	.dataa(!\altera_reset_synchronizer_int_chain[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\altera_reset_synchronizer_int_chain[4]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \altera_reset_synchronizer_int_chain[4]~0 .extended_lut = "off";
defparam \altera_reset_synchronizer_int_chain[4]~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \altera_reset_synchronizer_int_chain[4]~0 .shared_arith = "off";

dffeas \altera_reset_synchronizer_int_chain[4] (
	.clk(clk_clk),
	.d(\altera_reset_synchronizer_int_chain[4]~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[4]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[4] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[4] .power_up = "low";

dffeas \r_sync_rst_chain[3] (
	.clk(clk_clk),
	.d(\altera_reset_synchronizer_int_chain[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\r_sync_rst_chain[3]~q ),
	.prn(vcc));
defparam \r_sync_rst_chain[3] .is_wysiwyg = "true";
defparam \r_sync_rst_chain[3] .power_up = "low";

cyclonev_lcell_comb \r_sync_rst_chain~1 (
	.dataa(!\altera_reset_synchronizer_int_chain[2]~q ),
	.datab(!\r_sync_rst_chain[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\r_sync_rst_chain~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \r_sync_rst_chain~1 .extended_lut = "off";
defparam \r_sync_rst_chain~1 .lut_mask = 64'h7777777777777777;
defparam \r_sync_rst_chain~1 .shared_arith = "off";

dffeas \r_sync_rst_chain[2] (
	.clk(clk_clk),
	.d(\r_sync_rst_chain~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\r_sync_rst_chain[2]~q ),
	.prn(vcc));
defparam \r_sync_rst_chain[2] .is_wysiwyg = "true";
defparam \r_sync_rst_chain[2] .power_up = "low";

cyclonev_lcell_comb \r_sync_rst_chain~0 (
	.dataa(!\altera_reset_synchronizer_int_chain[2]~q ),
	.datab(!\r_sync_rst_chain[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\r_sync_rst_chain~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \r_sync_rst_chain~0 .extended_lut = "off";
defparam \r_sync_rst_chain~0 .lut_mask = 64'h7777777777777777;
defparam \r_sync_rst_chain~0 .shared_arith = "off";

dffeas \r_sync_rst_chain[1] (
	.clk(clk_clk),
	.d(\r_sync_rst_chain~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\r_sync_rst_chain[1]~q ),
	.prn(vcc));
defparam \r_sync_rst_chain[1] .is_wysiwyg = "true";
defparam \r_sync_rst_chain[1] .power_up = "low";

cyclonev_lcell_comb \WideOr0~0 (
	.dataa(!r_sync_rst1),
	.datab(!\altera_reset_synchronizer_int_chain[4]~q ),
	.datac(!\r_sync_rst_chain[1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr0~0 .extended_lut = "off";
defparam \WideOr0~0 .lut_mask = 64'hF7F7F7F7F7F7F7F7;
defparam \WideOr0~0 .shared_arith = "off";

cyclonev_lcell_comb \always2~0 (
	.dataa(!\r_sync_rst_chain[2]~q ),
	.datab(!\alt_rst_req_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always2~0 .extended_lut = "off";
defparam \always2~0 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \always2~0 .shared_arith = "off";

endmodule

module processor_altera_reset_synchronizer (
	altera_reset_synchronizer_int_chain_out1,
	altera_reset_synchronizer_int_chain_1,
	clk)/* synthesis synthesis_greybox=1 */;
output 	altera_reset_synchronizer_int_chain_out1;
output 	altera_reset_synchronizer_int_chain_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \altera_reset_synchronizer_int_chain[1]~q ;
wire \altera_reset_synchronizer_int_chain[0]~q ;


dffeas altera_reset_synchronizer_int_chain_out(
	.clk(clk),
	.d(\altera_reset_synchronizer_int_chain[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(altera_reset_synchronizer_int_chain_out1),
	.prn(vcc));
defparam altera_reset_synchronizer_int_chain_out.is_wysiwyg = "true";
defparam altera_reset_synchronizer_int_chain_out.power_up = "low";

cyclonev_lcell_comb \altera_reset_synchronizer_int_chain[1]~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(altera_reset_synchronizer_int_chain_1),
	.sumout(),
	.cout(),
	.shareout());
defparam \altera_reset_synchronizer_int_chain[1]~0 .extended_lut = "off";
defparam \altera_reset_synchronizer_int_chain[1]~0 .lut_mask = 64'h0000000000000000;
defparam \altera_reset_synchronizer_int_chain[1]~0 .shared_arith = "off";

dffeas \altera_reset_synchronizer_int_chain[1] (
	.clk(clk),
	.d(altera_reset_synchronizer_int_chain_1),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[1]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[1] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[1] .power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[0] (
	.clk(clk),
	.d(\altera_reset_synchronizer_int_chain[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[0]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[0] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[0] .power_up = "low";

endmodule

module processor_altera_reset_synchronizer_1 (
	altera_reset_synchronizer_int_chain_out1,
	clk,
	reset_reset_n)/* synthesis synthesis_greybox=1 */;
output 	altera_reset_synchronizer_int_chain_out1;
input 	clk;
input 	reset_reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \altera_reset_synchronizer_int_chain[1]~q ;
wire \altera_reset_synchronizer_int_chain[0]~q ;


dffeas altera_reset_synchronizer_int_chain_out(
	.clk(clk),
	.d(\altera_reset_synchronizer_int_chain[0]~q ),
	.asdata(vcc),
	.clrn(reset_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(altera_reset_synchronizer_int_chain_out1),
	.prn(vcc));
defparam altera_reset_synchronizer_int_chain_out.is_wysiwyg = "true";
defparam altera_reset_synchronizer_int_chain_out.power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[1] (
	.clk(clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(reset_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[1]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[1] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[1] .power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[0] (
	.clk(clk),
	.d(\altera_reset_synchronizer_int_chain[1]~q ),
	.asdata(vcc),
	.clrn(reset_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[0]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[0] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[0] .power_up = "low";

endmodule

module processor_processor_cpu (
	M_st_data_8,
	M_st_data_9,
	readdata_0,
	readdata_16,
	M_st_data_16,
	readdata_8,
	readdata_24,
	readdata_5,
	readdata_21,
	M_st_data_21,
	readdata_13,
	M_st_data_13,
	readdata_29,
	readdata_4,
	readdata_20,
	M_st_data_20,
	readdata_12,
	M_st_data_12,
	readdata_28,
	readdata_6,
	readdata_22,
	M_st_data_22,
	readdata_14,
	M_st_data_14,
	readdata_30,
	readdata_7,
	readdata_23,
	M_st_data_23,
	readdata_15,
	M_st_data_15,
	readdata_31,
	readdata_11,
	M_st_data_11,
	readdata_27,
	readdata_10,
	M_st_data_10,
	readdata_26,
	readdata_25,
	readdata_9,
	readdata_3,
	readdata_19,
	M_st_data_19,
	readdata_2,
	readdata_18,
	M_st_data_18,
	readdata_1,
	readdata_17,
	M_st_data_17,
	sr_0,
	ir_out_0,
	ir_out_1,
	M_st_data_0,
	r_sync_rst,
	clr_break_line1,
	d_write1,
	M_alu_result_5,
	M_alu_result_4,
	M_alu_result_6,
	M_alu_result_16,
	M_alu_result_15,
	M_alu_result_14,
	M_alu_result_13,
	M_alu_result_12,
	M_alu_result_11,
	M_alu_result_10,
	M_alu_result_9,
	M_alu_result_8,
	M_alu_result_7,
	M_alu_result_3,
	M_alu_result_2,
	M_st_data_1,
	M_st_data_2,
	M_st_data_3,
	M_st_data_4,
	M_st_data_5,
	M_st_data_6,
	M_st_data_7,
	d_read1,
	WideOr1,
	saved_grant_0,
	jtag_debug_module_waitrequest,
	mem_used_1,
	read_accepted,
	hbreak_enabled1,
	src2_valid,
	saved_grant_1,
	i_read1,
	has_pending_responses,
	ic_fill_tag_5,
	ic_fill_tag_4,
	ic_fill_tag_3,
	ic_fill_tag_2,
	ic_fill_tag_1,
	ic_fill_tag_0,
	Equal1,
	src0_valid,
	rf_source_valid,
	last_dest_id_1,
	d_readdata,
	WideOr0,
	nonposted_cmd_accepted,
	ic_fill_line_5,
	src_data_46,
	av_readdata_9,
	av_readdata_8,
	r_early_rst,
	timeout_occurred,
	control_register_0,
	ic_fill_line_0,
	ic_fill_line_1,
	ic_fill_line_2,
	ic_fill_line_3,
	ic_fill_line_4,
	ic_fill_ap_offset_0,
	ic_fill_ap_offset_1,
	ic_fill_ap_offset_2,
	M_mem_byte_en_0,
	M_mem_byte_en_2,
	M_mem_byte_en_1,
	M_st_data_24,
	M_mem_byte_en_3,
	src_payload,
	src_data_38,
	src_data_41,
	src_data_40,
	src_data_39,
	src_data_45,
	src_data_44,
	src_data_43,
	src_data_42,
	src_payload1,
	M_st_data_29,
	M_st_data_28,
	M_st_data_30,
	M_st_data_31,
	M_st_data_27,
	M_st_data_26,
	M_st_data_25,
	src_payload2,
	src_data_32,
	WideOr11,
	i_readdata,
	src_payload3,
	src_payload4,
	src_payload5,
	src_data_34,
	src_payload6,
	src_data_33,
	src_payload7,
	src_data_35,
	src_payload8,
	src_payload9,
	src_payload10,
	src_payload11,
	src_payload12,
	src_payload13,
	src_payload14,
	src_payload15,
	src_payload16,
	src_payload17,
	src_payload18,
	src_payload19,
	src_payload20,
	src_payload21,
	src_payload22,
	src_payload23,
	src_payload24,
	src_payload25,
	src_payload26,
	src_payload27,
	src_payload28,
	src_payload29,
	src_payload30,
	src_payload31,
	src_payload32,
	altera_internal_jtag,
	altera_internal_jtag1,
	state_1,
	state_4,
	virtual_ir_scan_reg,
	state_3,
	state_8,
	splitter_nodes_receive_1_3,
	irf_reg_0_2,
	irf_reg_1_2,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	M_st_data_8;
output 	M_st_data_9;
output 	readdata_0;
output 	readdata_16;
output 	M_st_data_16;
output 	readdata_8;
output 	readdata_24;
output 	readdata_5;
output 	readdata_21;
output 	M_st_data_21;
output 	readdata_13;
output 	M_st_data_13;
output 	readdata_29;
output 	readdata_4;
output 	readdata_20;
output 	M_st_data_20;
output 	readdata_12;
output 	M_st_data_12;
output 	readdata_28;
output 	readdata_6;
output 	readdata_22;
output 	M_st_data_22;
output 	readdata_14;
output 	M_st_data_14;
output 	readdata_30;
output 	readdata_7;
output 	readdata_23;
output 	M_st_data_23;
output 	readdata_15;
output 	M_st_data_15;
output 	readdata_31;
output 	readdata_11;
output 	M_st_data_11;
output 	readdata_27;
output 	readdata_10;
output 	M_st_data_10;
output 	readdata_26;
output 	readdata_25;
output 	readdata_9;
output 	readdata_3;
output 	readdata_19;
output 	M_st_data_19;
output 	readdata_2;
output 	readdata_18;
output 	M_st_data_18;
output 	readdata_1;
output 	readdata_17;
output 	M_st_data_17;
output 	sr_0;
output 	ir_out_0;
output 	ir_out_1;
output 	M_st_data_0;
input 	r_sync_rst;
output 	clr_break_line1;
output 	d_write1;
output 	M_alu_result_5;
output 	M_alu_result_4;
output 	M_alu_result_6;
output 	M_alu_result_16;
output 	M_alu_result_15;
output 	M_alu_result_14;
output 	M_alu_result_13;
output 	M_alu_result_12;
output 	M_alu_result_11;
output 	M_alu_result_10;
output 	M_alu_result_9;
output 	M_alu_result_8;
output 	M_alu_result_7;
output 	M_alu_result_3;
output 	M_alu_result_2;
output 	M_st_data_1;
output 	M_st_data_2;
output 	M_st_data_3;
output 	M_st_data_4;
output 	M_st_data_5;
output 	M_st_data_6;
output 	M_st_data_7;
output 	d_read1;
input 	WideOr1;
input 	saved_grant_0;
output 	jtag_debug_module_waitrequest;
input 	mem_used_1;
input 	read_accepted;
output 	hbreak_enabled1;
input 	src2_valid;
input 	saved_grant_1;
output 	i_read1;
input 	has_pending_responses;
output 	ic_fill_tag_5;
output 	ic_fill_tag_4;
output 	ic_fill_tag_3;
output 	ic_fill_tag_2;
output 	ic_fill_tag_1;
output 	ic_fill_tag_0;
input 	Equal1;
input 	src0_valid;
input 	rf_source_valid;
input 	last_dest_id_1;
input 	[31:0] d_readdata;
input 	WideOr0;
input 	nonposted_cmd_accepted;
output 	ic_fill_line_5;
input 	src_data_46;
input 	av_readdata_9;
input 	av_readdata_8;
input 	r_early_rst;
input 	timeout_occurred;
input 	control_register_0;
output 	ic_fill_line_0;
output 	ic_fill_line_1;
output 	ic_fill_line_2;
output 	ic_fill_line_3;
output 	ic_fill_line_4;
output 	ic_fill_ap_offset_0;
output 	ic_fill_ap_offset_1;
output 	ic_fill_ap_offset_2;
output 	M_mem_byte_en_0;
output 	M_mem_byte_en_2;
output 	M_mem_byte_en_1;
output 	M_st_data_24;
output 	M_mem_byte_en_3;
input 	src_payload;
input 	src_data_38;
input 	src_data_41;
input 	src_data_40;
input 	src_data_39;
input 	src_data_45;
input 	src_data_44;
input 	src_data_43;
input 	src_data_42;
input 	src_payload1;
output 	M_st_data_29;
output 	M_st_data_28;
output 	M_st_data_30;
output 	M_st_data_31;
output 	M_st_data_27;
output 	M_st_data_26;
output 	M_st_data_25;
input 	src_payload2;
input 	src_data_32;
input 	WideOr11;
input 	[31:0] i_readdata;
input 	src_payload3;
input 	src_payload4;
input 	src_payload5;
input 	src_data_34;
input 	src_payload6;
input 	src_data_33;
input 	src_payload7;
input 	src_data_35;
input 	src_payload8;
input 	src_payload9;
input 	src_payload10;
input 	src_payload11;
input 	src_payload12;
input 	src_payload13;
input 	src_payload14;
input 	src_payload15;
input 	src_payload16;
input 	src_payload17;
input 	src_payload18;
input 	src_payload19;
input 	src_payload20;
input 	src_payload21;
input 	src_payload22;
input 	src_payload23;
input 	src_payload24;
input 	src_payload25;
input 	src_payload26;
input 	src_payload27;
input 	src_payload28;
input 	src_payload29;
input 	src_payload30;
input 	src_payload31;
input 	src_payload32;
input 	altera_internal_jtag;
input 	altera_internal_jtag1;
input 	state_1;
input 	state_4;
input 	virtual_ir_scan_reg;
input 	state_3;
input 	state_8;
input 	splitter_nodes_receive_1_3;
input 	irf_reg_0_2;
input 	irf_reg_1_2;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \processor_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[0] ;
wire \processor_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[5] ;
wire \processor_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[5] ;
wire \processor_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[4] ;
wire \processor_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[4] ;
wire \processor_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[6] ;
wire \processor_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[6] ;
wire \processor_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[16] ;
wire \processor_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[16] ;
wire \processor_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[15] ;
wire \processor_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[15] ;
wire \processor_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[14] ;
wire \processor_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[14] ;
wire \processor_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[13] ;
wire \processor_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[13] ;
wire \processor_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[12] ;
wire \processor_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[12] ;
wire \processor_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[11] ;
wire \processor_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[11] ;
wire \processor_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[10] ;
wire \processor_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[10] ;
wire \processor_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[9] ;
wire \processor_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[9] ;
wire \processor_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[8] ;
wire \processor_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[8] ;
wire \processor_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[7] ;
wire \processor_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[7] ;
wire \processor_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[3] ;
wire \processor_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[3] ;
wire \processor_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[2] ;
wire \processor_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[2] ;
wire \processor_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[1] ;
wire \processor_cpu_ic_data|the_altsyncram|auto_generated|q_b[24] ;
wire \processor_cpu_ic_data|the_altsyncram|auto_generated|q_b[0] ;
wire \processor_cpu_ic_data|the_altsyncram|auto_generated|q_b[1] ;
wire \processor_cpu_ic_data|the_altsyncram|auto_generated|q_b[2] ;
wire \processor_cpu_ic_data|the_altsyncram|auto_generated|q_b[3] ;
wire \processor_cpu_ic_data|the_altsyncram|auto_generated|q_b[4] ;
wire \processor_cpu_ic_data|the_altsyncram|auto_generated|q_b[5] ;
wire \processor_cpu_ic_data|the_altsyncram|auto_generated|q_b[22] ;
wire \processor_cpu_ic_data|the_altsyncram|auto_generated|q_b[23] ;
wire \processor_cpu_ic_data|the_altsyncram|auto_generated|q_b[25] ;
wire \processor_cpu_ic_data|the_altsyncram|auto_generated|q_b[26] ;
wire \processor_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[0] ;
wire \processor_cpu_ic_data|the_altsyncram|auto_generated|q_b[14] ;
wire \processor_cpu_ic_tag|the_altsyncram|auto_generated|q_b[5] ;
wire \processor_cpu_ic_tag|the_altsyncram|auto_generated|q_b[1] ;
wire \processor_cpu_ic_tag|the_altsyncram|auto_generated|q_b[4] ;
wire \processor_cpu_ic_tag|the_altsyncram|auto_generated|q_b[0] ;
wire \processor_cpu_ic_tag|the_altsyncram|auto_generated|q_b[2] ;
wire \processor_cpu_ic_tag|the_altsyncram|auto_generated|q_b[3] ;
wire \processor_cpu_ic_data|the_altsyncram|auto_generated|q_b[12] ;
wire \processor_cpu_ic_data|the_altsyncram|auto_generated|q_b[11] ;
wire \processor_cpu_ic_data|the_altsyncram|auto_generated|q_b[16] ;
wire \processor_cpu_ic_data|the_altsyncram|auto_generated|q_b[15] ;
wire \processor_cpu_ic_data|the_altsyncram|auto_generated|q_b[13] ;
wire \processor_cpu_ic_data|the_altsyncram|auto_generated|q_b[21] ;
wire \processor_cpu_ic_data|the_altsyncram|auto_generated|q_b[29] ;
wire \processor_cpu_ic_data|the_altsyncram|auto_generated|q_b[27] ;
wire \processor_cpu_ic_data|the_altsyncram|auto_generated|q_b[28] ;
wire \processor_cpu_ic_data|the_altsyncram|auto_generated|q_b[30] ;
wire \processor_cpu_ic_data|the_altsyncram|auto_generated|q_b[31] ;
wire \processor_cpu_ic_data|the_altsyncram|auto_generated|q_b[10] ;
wire \processor_cpu_ic_data|the_altsyncram|auto_generated|q_b[6] ;
wire \processor_cpu_ic_data|the_altsyncram|auto_generated|q_b[8] ;
wire \processor_cpu_ic_data|the_altsyncram|auto_generated|q_b[7] ;
wire \processor_cpu_ic_data|the_altsyncram|auto_generated|q_b[20] ;
wire \processor_cpu_ic_data|the_altsyncram|auto_generated|q_b[19] ;
wire \processor_cpu_ic_data|the_altsyncram|auto_generated|q_b[18] ;
wire \processor_cpu_ic_data|the_altsyncram|auto_generated|q_b[17] ;
wire \processor_cpu_ic_data|the_altsyncram|auto_generated|q_b[9] ;
wire \processor_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[1] ;
wire \processor_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[31] ;
wire \processor_cpu_ic_tag|the_altsyncram|auto_generated|q_b[11] ;
wire \processor_cpu_ic_tag|the_altsyncram|auto_generated|q_b[13] ;
wire \processor_cpu_ic_tag|the_altsyncram|auto_generated|q_b[10] ;
wire \processor_cpu_ic_tag|the_altsyncram|auto_generated|q_b[12] ;
wire \ic_tag_wraddress[0]~q ;
wire \processor_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[17] ;
wire \processor_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[30] ;
wire \processor_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[31] ;
wire \ic_fill_valid_bits[5]~q ;
wire \ic_fill_valid_bits[7]~q ;
wire \ic_fill_valid_bits[4]~q ;
wire \processor_cpu_ic_tag|the_altsyncram|auto_generated|q_b[7] ;
wire \processor_cpu_ic_tag|the_altsyncram|auto_generated|q_b[9] ;
wire \processor_cpu_ic_tag|the_altsyncram|auto_generated|q_b[6] ;
wire \processor_cpu_ic_tag|the_altsyncram|auto_generated|q_b[8] ;
wire \ic_fill_valid_bits[6]~q ;
wire \processor_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[18] ;
wire \processor_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[17] ;
wire \processor_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[30] ;
wire \processor_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[29] ;
wire \processor_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[24] ;
wire \ic_fill_valid_bits[1]~q ;
wire \ic_fill_valid_bits[3]~q ;
wire \ic_fill_valid_bits[0]~q ;
wire \ic_fill_valid_bits[2]~q ;
wire \processor_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[21] ;
wire \processor_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[29] ;
wire \processor_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[20] ;
wire \processor_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[28] ;
wire \processor_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[22] ;
wire \processor_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[19] ;
wire \processor_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[18] ;
wire \processor_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[23] ;
wire \processor_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[27] ;
wire \processor_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[26] ;
wire \processor_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[25] ;
wire \processor_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[19] ;
wire \processor_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[28] ;
wire \processor_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[24] ;
wire \processor_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[21] ;
wire \processor_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[20] ;
wire \processor_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[22] ;
wire \processor_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[23] ;
wire \processor_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[27] ;
wire \processor_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[26] ;
wire \processor_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[25] ;
wire \the_processor_cpu_nios2_oci|the_processor_cpu_nios2_oci_debug|jtag_break~q ;
wire \the_processor_cpu_nios2_oci|the_processor_cpu_nios2_avalon_reg|oci_single_step_mode~q ;
wire \the_processor_cpu_nios2_oci|the_processor_cpu_nios2_avalon_reg|oci_ienable[16]~q ;
wire \the_processor_cpu_nios2_oci|the_processor_cpu_nios2_avalon_reg|oci_ienable[1]~q ;
wire \i_readdata_d1[24]~q ;
wire \i_readdata_d1[0]~q ;
wire \i_readdata_d1[1]~q ;
wire \i_readdata_d1[2]~q ;
wire \i_readdata_d1[3]~q ;
wire \i_readdata_d1[4]~q ;
wire \i_readdata_d1[5]~q ;
wire \i_readdata_d1[22]~q ;
wire \i_readdata_d1[23]~q ;
wire \i_readdata_d1[25]~q ;
wire \i_readdata_d1[26]~q ;
wire \i_readdata_d1[14]~q ;
wire \ic_tag_clr_valid_bits~q ;
wire \ic_tag_wren~combout ;
wire \ic_tag_wraddress[1]~q ;
wire \ic_tag_wraddress[2]~q ;
wire \ic_tag_wraddress[3]~q ;
wire \ic_tag_wraddress[4]~q ;
wire \ic_tag_wraddress[5]~q ;
wire \i_readdata_d1[12]~q ;
wire \i_readdata_d1[11]~q ;
wire \i_readdata_d1[16]~q ;
wire \i_readdata_d1[15]~q ;
wire \i_readdata_d1[13]~q ;
wire \i_readdata_d1[21]~q ;
wire \i_readdata_d1[29]~q ;
wire \i_readdata_d1[27]~q ;
wire \i_readdata_d1[28]~q ;
wire \i_readdata_d1[30]~q ;
wire \i_readdata_d1[31]~q ;
wire \i_readdata_d1[10]~q ;
wire \i_readdata_d1[6]~q ;
wire \i_readdata_d1[8]~q ;
wire \i_readdata_d1[7]~q ;
wire \i_readdata_d1[20]~q ;
wire \i_readdata_d1[19]~q ;
wire \i_readdata_d1[18]~q ;
wire \i_readdata_d1[17]~q ;
wire \i_readdata_d1[9]~q ;
wire \ic_tag_clr_valid_bits_nxt~combout ;
wire \ic_tag_wraddress_nxt~6_combout ;
wire \ic_tag_wraddress_nxt[1]~7_combout ;
wire \ic_tag_wraddress_nxt[1]~8_combout ;
wire \ic_tag_wraddress_nxt[2]~9_combout ;
wire \ic_tag_wraddress_nxt[3]~10_combout ;
wire \ic_tag_wraddress_nxt[4]~11_combout ;
wire \ic_tag_wraddress_nxt[5]~12_combout ;
wire \ic_fill_valid_bits_nxt~0_combout ;
wire \ic_fill_valid_bits_en~combout ;
wire \ic_fill_valid_bits_nxt~1_combout ;
wire \ic_fill_valid_bits_nxt~2_combout ;
wire \ic_fill_valid_bits_nxt~3_combout ;
wire \ic_fill_valid_bits_nxt~4_combout ;
wire \ic_fill_valid_bits_nxt~5_combout ;
wire \ic_fill_valid_bits_nxt~6_combout ;
wire \ic_fill_valid_bits_nxt~7_combout ;
wire \ic_tag_clr_valid_bits~0_combout ;
wire \F_iw[0]~2_combout ;
wire \F_iw[14]~12_combout ;
wire \av_ld_data_transfer~0_combout ;
wire \av_ld_aligning_data~q ;
wire \av_ld_or_div_done~q ;
wire \F_iw[5]~7_combout ;
wire \D_iw[5]~q ;
wire \E_iw[5]~q ;
wire \F_iw[4]~6_combout ;
wire \D_iw[4]~q ;
wire \E_iw[4]~q ;
wire \F_iw[3]~5_combout ;
wire \D_iw[3]~q ;
wire \E_iw[3]~q ;
wire \F_iw[2]~4_combout ;
wire \D_iw[2]~q ;
wire \E_iw[2]~q ;
wire \F_iw[1]~3_combout ;
wire \D_iw[1]~q ;
wire \E_iw[1]~q ;
wire \E_iw[0]~q ;
wire \Equal130~0_combout ;
wire \F_iw[12]~13_combout ;
wire \D_iw[12]~q ;
wire \E_iw[12]~q ;
wire \F_iw[11]~14_combout ;
wire \D_iw[11]~q ;
wire \E_iw[11]~q ;
wire \E_op_eret~0_combout ;
wire \F_iw[16]~15_combout ;
wire \D_iw[16]~q ;
wire \E_iw[16]~q ;
wire \F_iw[15]~16_combout ;
wire \D_iw[15]~q ;
wire \E_iw[15]~q ;
wire \F_iw[13]~17_combout ;
wire \D_iw[13]~q ;
wire \E_iw[13]~q ;
wire \E_hbreak_req~0_combout ;
wire \wait_for_one_post_bret_inst~0_combout ;
wire \wait_for_one_post_bret_inst~q ;
wire \hbreak_req~0_combout ;
wire \E_valid~1_combout ;
wire \M_valid_from_E~q ;
wire \D_ctrl_ld~0_combout ;
wire \E_ctrl_ld~q ;
wire \M_ctrl_ld~q ;
wire \M_status_reg_pie~0_combout ;
wire \Equal4~0_combout ;
wire \D_ctrl_shift_logical~0_combout ;
wire \E_ctrl_shift_rot~q ;
wire \D_ctrl_b_not_src~0_combout ;
wire \D_wr_dst_reg~1_combout ;
wire \D_ctrl_src2_choose_imm~combout ;
wire \E_ctrl_src2_choose_imm~q ;
wire \F_iw[6]~25_combout ;
wire \D_iw[6]~q ;
wire \D_ctrl_hi_imm16~0_combout ;
wire \E_src2_imm[0]~q ;
wire \M_ctrl_shift_rot~q ;
wire \d_readdata_d1[3]~q ;
wire \d_readdata_d1[19]~q ;
wire \d_readdata_d1[11]~q ;
wire \d_readdata_d1[27]~q ;
wire \D_ctrl_crst~0_combout ;
wire \Equal107~1_combout ;
wire \E_ctrl_rdctl_inst~q ;
wire \D_ctrl_implicit_dst_retaddr~0_combout ;
wire \D_ctrl_retaddr~0_combout ;
wire \D_ctrl_break~0_combout ;
wire \Equal4~1_combout ;
wire \Equal107~0_combout ;
wire \D_ctrl_implicit_dst_eretaddr~0_combout ;
wire \D_ctrl_exception~0_combout ;
wire \D_ctrl_retaddr~1_combout ;
wire \E_ctrl_retaddr~q ;
wire \Equal4~5_combout ;
wire \Equal4~6_combout ;
wire \Equal4~7_combout ;
wire \Equal4~8_combout ;
wire \Equal4~9_combout ;
wire \Equal4~10_combout ;
wire \D_ctrl_cmp~0_combout ;
wire \D_ctrl_cmp~1_combout ;
wire \D_ctrl_cmp~2_combout ;
wire \E_ctrl_cmp~q ;
wire \E_alu_result~0_combout ;
wire \D_ctrl_alu_subtract~0_combout ;
wire \D_ctrl_alu_subtract~1_combout ;
wire \E_ctrl_alu_subtract~q ;
wire \d_readdata_d1[1]~q ;
wire \d_readdata_d1[17]~q ;
wire \d_readdata_d1[9]~q ;
wire \d_readdata_d1[25]~q ;
wire \D_compare_op[1]~0_combout ;
wire \E_compare_op[1]~q ;
wire \D_compare_op[0]~1_combout ;
wire \E_compare_op[0]~q ;
wire \D_ctrl_a_not_src~0_combout ;
wire \F_iw[29]~19_combout ;
wire \D_iw[29]~q ;
wire \F_iw[23]~9_combout ;
wire \D_iw[23]~q ;
wire \F_iw[18]~30_combout ;
wire \D_iw[18]~q ;
wire \D_ctrl_implicit_dst_eretaddr~1_combout ;
wire \D_ctrl_implicit_dst_eretaddr~2_combout ;
wire \D_dst_regnum[1]~2_combout ;
wire \F_iw[22]~8_combout ;
wire \D_iw[22]~q ;
wire \F_iw[17]~31_combout ;
wire \D_iw[17]~q ;
wire \D_dst_regnum[4]~0_combout ;
wire \D_dst_regnum[0]~3_combout ;
wire \F_iw[25]~10_combout ;
wire \D_iw[25]~q ;
wire \F_iw[20]~28_combout ;
wire \D_iw[20]~q ;
wire \D_dst_regnum[3]~4_combout ;
wire \F_iw[26]~11_combout ;
wire \D_iw[26]~q ;
wire \F_iw[21]~18_combout ;
wire \D_iw[21]~q ;
wire \D_dst_regnum[4]~5_combout ;
wire \D_wr_dst_reg~0_combout ;
wire \D_wr_dst_reg~combout ;
wire \E_wr_dst_reg_from_D~q ;
wire \E_wr_dst_reg~0_combout ;
wire \E_dst_regnum[0]~q ;
wire \E_dst_regnum[1]~q ;
wire \F_iw[27]~20_combout ;
wire \D_iw[27]~q ;
wire \F_iw[28]~21_combout ;
wire \D_iw[28]~q ;
wire \D_src1_hazard_E~0_combout ;
wire \E_dst_regnum[3]~q ;
wire \E_dst_regnum[4]~q ;
wire \F_iw[30]~22_combout ;
wire \D_iw[30]~q ;
wire \F_iw[31]~23_combout ;
wire \D_iw[31]~q ;
wire \D_src1_hazard_E~1_combout ;
wire \D_src1_hazard_E~combout ;
wire \E_src1_hazard_M~q ;
wire \D_ctrl_shift_rot_right~0_combout ;
wire \E_ctrl_shift_rot_right~q ;
wire \M_ctrl_shift_rot_right~q ;
wire \D_ctrl_shift_logical~1_combout ;
wire \E_ctrl_shift_logical~q ;
wire \M_ctrl_shift_logical~q ;
wire \D_ctrl_rot_right~0_combout ;
wire \E_ctrl_rot_right~q ;
wire \M_ctrl_rot_right~q ;
wire \M_shift_rot_fill_bit~0_combout ;
wire \d_readdata_d1[31]~q ;
wire \d_readdata_d1[15]~q ;
wire \d_readdata_d1[23]~q ;
wire \M_iw[4]~q ;
wire \M_iw[3]~q ;
wire \av_sign_bit~0_combout ;
wire \D_ctrl_b_is_dst~0_combout ;
wire \E_ctrl_ld_signed~q ;
wire \M_ctrl_ld_signed~q ;
wire \d_readdata_d1[7]~q ;
wire \av_fill_bit~0_combout ;
wire \d_readdata_d1[30]~q ;
wire \av_ld_data_aligned_or_div[30]~q ;
wire \E_stw_data[30]~15_combout ;
wire \M_wr_data_unfiltered[30]~19_combout ;
wire \M_dst_regnum[4]~q ;
wire \M_wr_dst_reg~q ;
wire \M_dst_regnum[0]~q ;
wire \M_dst_regnum[1]~q ;
wire \D_src2_hazard_M~0_combout ;
wire \M_dst_regnum[2]~q ;
wire \M_dst_regnum[3]~q ;
wire \D_src2_hazard_M~1_combout ;
wire \D_src2_hazard_M~combout ;
wire \W_dst_regnum[4]~q ;
wire \W_wr_dst_reg~0_combout ;
wire \W_wr_dst_reg~q ;
wire \W_dst_regnum[0]~q ;
wire \W_dst_regnum[1]~q ;
wire \D_src2_hazard_W~0_combout ;
wire \W_dst_regnum[2]~q ;
wire \W_dst_regnum[3]~q ;
wire \D_src2_hazard_W~1_combout ;
wire \D_src2_hazard_W~combout ;
wire \W_wr_data[30]~q ;
wire \D_src2_prelim[30]~19_combout ;
wire \E_src2_prelim[30]~q ;
wire \E_stw_data[30]~16_combout ;
wire \E_stw_data[30]~17_combout ;
wire \D_ctrl_logic~1_combout ;
wire \D_ctrl_unsigned_lo_imm16~combout ;
wire \Equal171~0_combout ;
wire \E_src2_imm[30]~q ;
wire \d_readdata_d1[28]~q ;
wire \av_ld_data_aligned_or_div[28]~q ;
wire \E_stw_data[28]~26_combout ;
wire \M_wr_data_unfiltered[28]~29_combout ;
wire \W_wr_data[28]~q ;
wire \D_src2_prelim[28]~24_combout ;
wire \E_src2_prelim[28]~q ;
wire \E_stw_data[28]~27_combout ;
wire \E_stw_data[28]~28_combout ;
wire \E_src2_imm[28]~q ;
wire \d_readdata_d1[26]~q ;
wire \av_ld_data_aligned_or_div[26]~q ;
wire \E_stw_data[26]~38_combout ;
wire \M_wr_data_unfiltered[26]~31_combout ;
wire \W_wr_data[26]~q ;
wire \D_src2_prelim[26]~29_combout ;
wire \E_src2_prelim[26]~q ;
wire \E_stw_data[26]~39_combout ;
wire \E_stw_data[26]~40_combout ;
wire \E_src2_imm[26]~q ;
wire \d_readdata_d1[24]~q ;
wire \av_ld_data_aligned_or_div[24]~q ;
wire \E_stw_data[24]~18_combout ;
wire \M_wr_data_unfiltered[24]~27_combout ;
wire \W_wr_data[24]~q ;
wire \D_src2_prelim[24]~20_combout ;
wire \E_src2_prelim[24]~q ;
wire \E_stw_data[24]~19_combout ;
wire \E_stw_data[24]~20_combout ;
wire \E_src2_imm[24]~q ;
wire \d_readdata_d1[22]~q ;
wire \av_ld_data_aligned_or_div[22]~q ;
wire \E_stw_data[22]~29_combout ;
wire \M_wr_data_unfiltered[22]~30_combout ;
wire \W_wr_data[22]~q ;
wire \D_src2_prelim[22]~25_combout ;
wire \E_src2_prelim[22]~q ;
wire \E_stw_data[22]~30_combout ;
wire \E_stw_data[22]~31_combout ;
wire \E_src2_imm[22]~q ;
wire \d_readdata_d1[20]~q ;
wire \av_ld_data_aligned_or_div[20]~q ;
wire \E_stw_data[20]~23_combout ;
wire \M_wr_data_unfiltered[20]~28_combout ;
wire \W_wr_data[20]~q ;
wire \D_src2_prelim[20]~23_combout ;
wire \E_src2_prelim[20]~q ;
wire \E_stw_data[20]~24_combout ;
wire \E_stw_data[20]~25_combout ;
wire \F_iw[10]~24_combout ;
wire \D_iw[10]~q ;
wire \E_src2_imm[20]~q ;
wire \d_readdata_d1[18]~q ;
wire \av_ld_data_aligned_or_div[18]~q ;
wire \E_stw_data[18]~32_combout ;
wire \M_wr_data_unfiltered[18]~23_combout ;
wire \W_wr_data[18]~q ;
wire \D_src2_prelim[18]~26_combout ;
wire \E_src2_prelim[18]~q ;
wire \E_stw_data[18]~33_combout ;
wire \E_stw_data[18]~34_combout ;
wire \F_iw[8]~26_combout ;
wire \D_iw[8]~q ;
wire \E_src2_imm[18]~q ;
wire \d_readdata_d1[16]~q ;
wire \av_ld_data_aligned_or_div[16]~q ;
wire \E_src1[16]~7_combout ;
wire \M_wr_data_unfiltered[16]~13_combout ;
wire \D_src1_hazard_M~0_combout ;
wire \D_src1_hazard_M~1_combout ;
wire \D_src1_hazard_M~combout ;
wire \D_src1_hazard_W~0_combout ;
wire \D_src1_hazard_W~1_combout ;
wire \D_src1_hazard_W~combout ;
wire \W_wr_data[16]~q ;
wire \D_src1_prelim[16]~3_combout ;
wire \E_src1_prelim[16]~q ;
wire \E_src1[16]~8_combout ;
wire \E_src1[16]~9_combout ;
wire \Equal2~0_combout ;
wire \av_ld_byte1_data[7]~0_combout ;
wire \av_ld_data_aligned_or_div[15]~q ;
wire \M_wr_data_unfiltered[15]~1_combout ;
wire \W_wr_data[15]~q ;
wire \D_src1_prelim[15]~4_combout ;
wire \E_src1_prelim[15]~q ;
wire \E_src1[15]~10_combout ;
wire \d_readdata_d1[14]~q ;
wire \av_ld_byte1_data[6]~1_combout ;
wire \av_ld_data_aligned_or_div[14]~q ;
wire \M_wr_data_unfiltered[14]~2_combout ;
wire \W_wr_data[14]~q ;
wire \D_src1_prelim[14]~5_combout ;
wire \E_src1_prelim[14]~q ;
wire \E_src1[14]~11_combout ;
wire \d_readdata_d1[12]~q ;
wire \av_ld_byte1_data[4]~3_combout ;
wire \av_ld_data_aligned_or_div[12]~q ;
wire \M_wr_data_unfiltered[12]~4_combout ;
wire \W_wr_data[12]~q ;
wire \D_src1_prelim[12]~7_combout ;
wire \E_src1_prelim[12]~q ;
wire \E_src1[12]~13_combout ;
wire \av_ld_byte1_data[3]~4_combout ;
wire \av_ld_data_aligned_or_div[11]~q ;
wire \M_wr_data_unfiltered[11]~5_combout ;
wire \W_wr_data[11]~q ;
wire \D_src1_prelim[11]~8_combout ;
wire \E_src1_prelim[11]~q ;
wire \E_src1[11]~14_combout ;
wire \d_readdata_d1[10]~q ;
wire \av_ld_byte1_data[2]~5_combout ;
wire \av_ld_data_aligned_or_div[10]~q ;
wire \E_src1[10]~15_combout ;
wire \M_wr_data_unfiltered[10]~14_combout ;
wire \W_wr_data[10]~q ;
wire \D_src1_prelim[10]~9_combout ;
wire \E_src1_prelim[10]~q ;
wire \E_src1[10]~16_combout ;
wire \E_src1[10]~17_combout ;
wire \av_ld_byte1_data[1]~6_combout ;
wire \av_ld_data_aligned_or_div[9]~q ;
wire \M_wr_data_unfiltered[9]~6_combout ;
wire \W_wr_data[9]~q ;
wire \D_src1_prelim[9]~10_combout ;
wire \E_src1_prelim[9]~q ;
wire \E_src1[9]~18_combout ;
wire \d_readdata_d1[8]~q ;
wire \av_ld_byte1_data[0]~7_combout ;
wire \av_ld_data_aligned_or_div[8]~q ;
wire \E_src1[8]~19_combout ;
wire \M_wr_data_unfiltered[8]~15_combout ;
wire \W_wr_data[8]~q ;
wire \D_src1_prelim[8]~11_combout ;
wire \E_src1_prelim[8]~q ;
wire \E_src1[8]~20_combout ;
wire \E_src1[8]~21_combout ;
wire \d_readdata_d1[5]~q ;
wire \d_readdata_d1[21]~q ;
wire \d_readdata_d1[13]~q ;
wire \d_readdata_d1[29]~q ;
wire \av_ld_byte0_data[5]~1_combout ;
wire \av_ld_data_aligned_or_div[5]~q ;
wire \M_wr_data_unfiltered[5]~0_combout ;
wire \W_wr_data[5]~q ;
wire \D_src1_prelim[5]~0_combout ;
wire \E_src1_prelim[5]~q ;
wire \E_src1[5]~0_combout ;
wire \d_readdata_d1[4]~q ;
wire \av_ld_byte0_data[4]~2_combout ;
wire \av_ld_data_aligned_or_div[4]~q ;
wire \E_src1[4]~1_combout ;
wire \M_wr_data_unfiltered[4]~11_combout ;
wire \W_wr_data[4]~q ;
wire \D_src1_prelim[4]~1_combout ;
wire \E_src1_prelim[4]~q ;
wire \E_src1[4]~2_combout ;
wire \E_src1[4]~3_combout ;
wire \M_shift_rot_result_nxt[4]~2_combout ;
wire \M_shift_rot_result[4]~q ;
wire \M_shift_rot_result_nxt[5]~1_combout ;
wire \M_shift_rot_result[5]~q ;
wire \d_readdata_d1[6]~q ;
wire \av_ld_byte0_data[6]~3_combout ;
wire \av_ld_data_aligned_or_div[6]~q ;
wire \E_src1[6]~4_combout ;
wire \M_wr_data_unfiltered[6]~12_combout ;
wire \W_wr_data[6]~q ;
wire \D_src1_prelim[6]~2_combout ;
wire \E_src1_prelim[6]~q ;
wire \E_src1[6]~5_combout ;
wire \E_src1[6]~6_combout ;
wire \M_shift_rot_result_nxt[6]~3_combout ;
wire \M_shift_rot_result[6]~q ;
wire \av_ld_byte0_data[7]~4_combout ;
wire \av_ld_data_aligned_or_div[7]~q ;
wire \M_wr_data_unfiltered[7]~7_combout ;
wire \W_wr_data[7]~q ;
wire \D_src1_prelim[7]~12_combout ;
wire \E_src1_prelim[7]~q ;
wire \E_src1[7]~22_combout ;
wire \M_shift_rot_result_nxt[7]~13_combout ;
wire \M_shift_rot_result[7]~q ;
wire \M_shift_rot_result_nxt[8]~12_combout ;
wire \M_shift_rot_result[8]~q ;
wire \M_shift_rot_result_nxt[9]~11_combout ;
wire \M_shift_rot_result[9]~q ;
wire \M_shift_rot_result_nxt[10]~10_combout ;
wire \M_shift_rot_result[10]~q ;
wire \M_shift_rot_result_nxt[11]~9_combout ;
wire \M_shift_rot_result[11]~q ;
wire \M_shift_rot_result_nxt[12]~8_combout ;
wire \M_shift_rot_result[12]~q ;
wire \av_ld_byte1_data[5]~2_combout ;
wire \av_ld_data_aligned_or_div[13]~q ;
wire \M_wr_data_unfiltered[13]~3_combout ;
wire \W_wr_data[13]~q ;
wire \D_src1_prelim[13]~6_combout ;
wire \E_src1_prelim[13]~q ;
wire \E_src1[13]~12_combout ;
wire \M_shift_rot_result_nxt[13]~7_combout ;
wire \M_shift_rot_result[13]~q ;
wire \M_shift_rot_result_nxt[14]~6_combout ;
wire \M_shift_rot_result[14]~q ;
wire \M_shift_rot_result_nxt[15]~5_combout ;
wire \M_shift_rot_result[15]~q ;
wire \M_shift_rot_result_nxt[16]~4_combout ;
wire \M_shift_rot_result[16]~q ;
wire \W_wr_data[17]~q ;
wire \D_src1_prelim[17]~18_combout ;
wire \E_src1_prelim[17]~q ;
wire \E_src1[17]~32_combout ;
wire \M_shift_rot_result_nxt[17]~18_combout ;
wire \M_shift_rot_result[17]~q ;
wire \av_ld_data_aligned_or_div[17]~q ;
wire \F_iw[7]~27_combout ;
wire \D_iw[7]~q ;
wire \E_src2_imm[17]~q ;
wire \E_stw_data[16]~0_combout ;
wire \D_src2_prelim[16]~4_combout ;
wire \E_src2_prelim[16]~q ;
wire \E_stw_data[16]~1_combout ;
wire \E_stw_data[16]~2_combout ;
wire \E_src2_imm[16]~q ;
wire \D_src2_prelim[15]~5_combout ;
wire \E_src2_prelim[15]~q ;
wire \E_stw_data[15]~3_combout ;
wire \E_src2_imm[15]~q ;
wire \D_src2_prelim[14]~6_combout ;
wire \E_src2_prelim[14]~q ;
wire \E_stw_data[14]~4_combout ;
wire \E_src2_imm[14]~q ;
wire \D_src2_prelim[13]~7_combout ;
wire \E_src2_prelim[13]~q ;
wire \E_stw_data[13]~13_combout ;
wire \F_iw[19]~29_combout ;
wire \D_iw[19]~q ;
wire \E_src2_imm[13]~q ;
wire \D_src2_prelim[12]~8_combout ;
wire \E_src2_prelim[12]~q ;
wire \E_stw_data[12]~5_combout ;
wire \E_src2_imm[12]~q ;
wire \D_src2_prelim[11]~9_combout ;
wire \E_src2_prelim[11]~q ;
wire \E_stw_data[11]~14_combout ;
wire \E_src2_imm[11]~q ;
wire \E_stw_data[10]~6_combout ;
wire \D_src2_prelim[10]~10_combout ;
wire \E_src2_prelim[10]~q ;
wire \E_stw_data[10]~7_combout ;
wire \E_stw_data[10]~8_combout ;
wire \E_src2_imm[10]~q ;
wire \D_src2_prelim[9]~11_combout ;
wire \E_src2_prelim[9]~q ;
wire \E_stw_data[9]~12_combout ;
wire \E_src2_imm[9]~q ;
wire \E_stw_data[8]~9_combout ;
wire \D_src2_prelim[8]~12_combout ;
wire \E_src2_prelim[8]~q ;
wire \E_stw_data[8]~10_combout ;
wire \E_stw_data[8]~11_combout ;
wire \E_src2_imm[8]~q ;
wire \D_src2_prelim[7]~13_combout ;
wire \E_src2_prelim[7]~q ;
wire \E_stb_data[7]~15_combout ;
wire \E_src2_imm[7]~q ;
wire \E_stb_data[6]~6_combout ;
wire \D_src2_prelim[6]~3_combout ;
wire \E_src2_prelim[6]~q ;
wire \E_stb_data[6]~7_combout ;
wire \E_stb_data[6]~8_combout ;
wire \E_src2_imm[6]~q ;
wire \D_src2_prelim[5]~1_combout ;
wire \E_src2_prelim[5]~q ;
wire \E_stb_data[5]~14_combout ;
wire \E_src2_imm[5]~q ;
wire \E_stb_data[4]~3_combout ;
wire \D_src2_prelim[4]~2_combout ;
wire \E_src2_prelim[4]~q ;
wire \E_stb_data[4]~4_combout ;
wire \E_stb_data[4]~5_combout ;
wire \E_src2_imm[4]~q ;
wire \W_wr_data[3]~q ;
wire \D_src2_prelim[3]~14_combout ;
wire \E_src2_prelim[3]~q ;
wire \E_stb_data[3]~13_combout ;
wire \F_iw[9]~32_combout ;
wire \D_iw[9]~q ;
wire \E_src2_imm[3]~q ;
wire \d_readdata_d1[2]~q ;
wire \av_ld_byte0_data[2]~6_combout ;
wire \av_ld_data_aligned_or_div[2]~q ;
wire \E_stb_data[2]~9_combout ;
wire \M_wr_data_unfiltered[2]~16_combout ;
wire \W_wr_data[2]~q ;
wire \D_src2_prelim[2]~15_combout ;
wire \E_src2_prelim[2]~q ;
wire \E_stb_data[2]~10_combout ;
wire \E_stb_data[2]~11_combout ;
wire \E_src2_imm[2]~q ;
wire \E_src1[2]~24_combout ;
wire \D_src1_prelim[2]~14_combout ;
wire \E_src1_prelim[2]~q ;
wire \E_src1[2]~25_combout ;
wire \E_src1[2]~26_combout ;
wire \E_src2_imm[1]~q ;
wire \W_wr_data[1]~q ;
wire \D_src1_prelim[1]~16_combout ;
wire \E_src1_prelim[1]~q ;
wire \E_src1[1]~30_combout ;
wire \d_readdata_d1[0]~q ;
wire \av_ld_byte0_data[0]~0_combout ;
wire \av_ld_data_aligned_or_div[0]~q ;
wire \E_src1[0]~27_combout ;
wire \W_wr_data[0]~q ;
wire \D_src1_prelim[0]~15_combout ;
wire \E_src1_prelim[0]~q ;
wire \E_src1[0]~28_combout ;
wire \E_src1[0]~29_combout ;
wire \Add8~78_cout ;
wire \Add8~66 ;
wire \Add8~70 ;
wire \Add8~58 ;
wire \Add8~54 ;
wire \Add8~6 ;
wire \Add8~2 ;
wire \Add8~10 ;
wire \Add8~50 ;
wire \Add8~46 ;
wire \Add8~42 ;
wire \Add8~38 ;
wire \Add8~34 ;
wire \Add8~30 ;
wire \Add8~26 ;
wire \Add8~22 ;
wire \Add8~18 ;
wire \Add8~14 ;
wire \Add8~85_sumout ;
wire \D_src2_prelim[17]~18_combout ;
wire \E_src2_prelim[17]~q ;
wire \E_arith_src2[17]~13_combout ;
wire \E_alu_result[17]~28_combout ;
wire \E_alu_result[17]~29_combout ;
wire \M_alu_result[17]~q ;
wire \M_wr_data_unfiltered[17]~18_combout ;
wire \E_stw_data[17]~35_combout ;
wire \Add8~86 ;
wire \Add8~93_sumout ;
wire \E_alu_result[18]~32_combout ;
wire \E_alu_result[18]~33_combout ;
wire \M_alu_result[18]~q ;
wire \E_src1[18]~36_combout ;
wire \D_src1_prelim[18]~20_combout ;
wire \E_src1_prelim[18]~q ;
wire \E_src1[18]~37_combout ;
wire \E_src1[18]~38_combout ;
wire \M_shift_rot_result_nxt[18]~20_combout ;
wire \M_shift_rot_result[18]~q ;
wire \W_wr_data[19]~q ;
wire \D_src1_prelim[19]~22_combout ;
wire \E_src1_prelim[19]~q ;
wire \E_src1[19]~40_combout ;
wire \M_shift_rot_result_nxt[19]~22_combout ;
wire \M_shift_rot_result[19]~q ;
wire \av_ld_data_aligned_or_div[19]~q ;
wire \E_src2_imm[19]~q ;
wire \Add8~94 ;
wire \Add8~117_sumout ;
wire \D_src2_prelim[19]~31_combout ;
wire \E_src2_prelim[19]~q ;
wire \E_arith_src2[19]~16_combout ;
wire \E_alu_result[19]~46_combout ;
wire \E_alu_result[19]~47_combout ;
wire \M_alu_result[19]~q ;
wire \M_wr_data_unfiltered[19]~22_combout ;
wire \E_stw_data[19]~42_combout ;
wire \Add8~118 ;
wire \Add8~109_sumout ;
wire \E_alu_result[20]~40_combout ;
wire \E_alu_result[20]~41_combout ;
wire \M_alu_result[20]~q ;
wire \E_src1[20]~48_combout ;
wire \D_src1_prelim[20]~26_combout ;
wire \E_src1_prelim[20]~q ;
wire \E_src1[20]~49_combout ;
wire \E_src1[20]~50_combout ;
wire \M_shift_rot_result_nxt[20]~26_combout ;
wire \M_shift_rot_result[20]~q ;
wire \W_wr_data[21]~q ;
wire \D_src1_prelim[21]~25_combout ;
wire \E_src1_prelim[21]~q ;
wire \E_src1[21]~47_combout ;
wire \M_shift_rot_result_nxt[21]~25_combout ;
wire \M_shift_rot_result[21]~q ;
wire \av_ld_data_aligned_or_div[21]~q ;
wire \E_src2_imm[21]~q ;
wire \Add8~110 ;
wire \Add8~105_sumout ;
wire \D_src2_prelim[21]~21_combout ;
wire \E_src2_prelim[21]~q ;
wire \E_arith_src2[21]~15_combout ;
wire \E_alu_result[21]~38_combout ;
wire \E_alu_result[21]~39_combout ;
wire \M_alu_result[21]~q ;
wire \M_wr_data_unfiltered[21]~21_combout ;
wire \E_stw_data[21]~21_combout ;
wire \Add8~106 ;
wire \Add8~113_sumout ;
wire \E_alu_result[22]~44_combout ;
wire \E_alu_result[22]~45_combout ;
wire \M_alu_result[22]~q ;
wire \E_src1[22]~51_combout ;
wire \D_src1_prelim[22]~27_combout ;
wire \E_src1_prelim[22]~q ;
wire \E_src1[22]~52_combout ;
wire \E_src1[22]~53_combout ;
wire \M_shift_rot_result_nxt[22]~27_combout ;
wire \M_shift_rot_result[22]~q ;
wire \W_wr_data[23]~q ;
wire \D_src1_prelim[23]~28_combout ;
wire \E_src1_prelim[23]~q ;
wire \E_src1[23]~54_combout ;
wire \M_shift_rot_result_nxt[23]~28_combout ;
wire \M_shift_rot_result[23]~q ;
wire \av_ld_data_aligned_or_div[23]~q ;
wire \E_src2_imm[23]~q ;
wire \Add8~114 ;
wire \Add8~121_sumout ;
wire \D_src2_prelim[23]~27_combout ;
wire \E_src2_prelim[23]~q ;
wire \E_arith_src2[23]~17_combout ;
wire \E_alu_result[23]~48_combout ;
wire \E_alu_result[23]~49_combout ;
wire \M_alu_result[23]~q ;
wire \M_wr_data_unfiltered[23]~24_combout ;
wire \E_stw_data[23]~36_combout ;
wire \Add8~122 ;
wire \Add8~97_sumout ;
wire \E_alu_result[24]~36_combout ;
wire \E_alu_result[24]~37_combout ;
wire \M_alu_result[24]~q ;
wire \E_src1[24]~44_combout ;
wire \D_src1_prelim[24]~24_combout ;
wire \E_src1_prelim[24]~q ;
wire \E_src1[24]~45_combout ;
wire \E_src1[24]~46_combout ;
wire \M_shift_rot_result_nxt[24]~24_combout ;
wire \M_shift_rot_result[24]~q ;
wire \W_wr_data[25]~q ;
wire \D_src1_prelim[25]~31_combout ;
wire \E_src1_prelim[25]~q ;
wire \E_src1[25]~59_combout ;
wire \M_shift_rot_result_nxt[25]~31_combout ;
wire \M_shift_rot_result[25]~q ;
wire \av_ld_data_aligned_or_div[25]~q ;
wire \E_src2_imm[25]~q ;
wire \Add8~98 ;
wire \Add8~133_sumout ;
wire \D_src2_prelim[25]~30_combout ;
wire \E_src2_prelim[25]~q ;
wire \E_arith_src2[25]~19_combout ;
wire \E_alu_result[25]~54_combout ;
wire \E_alu_result[25]~55_combout ;
wire \M_alu_result[25]~q ;
wire \M_wr_data_unfiltered[25]~26_combout ;
wire \E_stw_data[25]~41_combout ;
wire \Add8~134 ;
wire \Add8~129_sumout ;
wire \E_alu_result[26]~52_combout ;
wire \E_alu_result[26]~53_combout ;
wire \M_alu_result[26]~q ;
wire \E_src1[26]~56_combout ;
wire \D_src1_prelim[26]~30_combout ;
wire \E_src1_prelim[26]~q ;
wire \E_src1[26]~57_combout ;
wire \E_src1[26]~58_combout ;
wire \M_shift_rot_result_nxt[26]~30_combout ;
wire \M_shift_rot_result[26]~q ;
wire \W_wr_data[27]~q ;
wire \D_src1_prelim[27]~29_combout ;
wire \E_src1_prelim[27]~q ;
wire \E_src1[27]~55_combout ;
wire \M_shift_rot_result_nxt[27]~29_combout ;
wire \M_shift_rot_result[27]~q ;
wire \av_ld_data_aligned_or_div[27]~q ;
wire \E_src2_imm[27]~q ;
wire \Add8~130 ;
wire \Add8~125_sumout ;
wire \D_src2_prelim[27]~28_combout ;
wire \E_src2_prelim[27]~q ;
wire \E_arith_src2[27]~18_combout ;
wire \E_alu_result[27]~50_combout ;
wire \E_alu_result[27]~51_combout ;
wire \M_alu_result[27]~q ;
wire \M_wr_data_unfiltered[27]~25_combout ;
wire \E_stw_data[27]~37_combout ;
wire \Add8~126 ;
wire \Add8~101_sumout ;
wire \E_alu_result[28]~42_combout ;
wire \E_alu_result[28]~43_combout ;
wire \M_alu_result[28]~q ;
wire \E_src1[28]~41_combout ;
wire \D_src1_prelim[28]~23_combout ;
wire \E_src1_prelim[28]~q ;
wire \E_src1[28]~42_combout ;
wire \E_src1[28]~43_combout ;
wire \M_shift_rot_result_nxt[28]~23_combout ;
wire \M_shift_rot_result[28]~q ;
wire \W_wr_data[29]~q ;
wire \D_src1_prelim[29]~21_combout ;
wire \E_src1_prelim[29]~q ;
wire \E_src1[29]~39_combout ;
wire \M_shift_rot_result_nxt[29]~21_combout ;
wire \M_shift_rot_result[29]~q ;
wire \av_ld_data_aligned_or_div[29]~q ;
wire \E_src2_imm[29]~q ;
wire \Add8~102 ;
wire \Add8~89_sumout ;
wire \D_src2_prelim[29]~22_combout ;
wire \E_src2_prelim[29]~q ;
wire \E_arith_src2[29]~14_combout ;
wire \E_alu_result[29]~34_combout ;
wire \E_alu_result[29]~35_combout ;
wire \M_alu_result[29]~q ;
wire \M_wr_data_unfiltered[29]~20_combout ;
wire \E_stw_data[29]~22_combout ;
wire \Add8~90 ;
wire \Add8~81_sumout ;
wire \E_alu_result[30]~30_combout ;
wire \E_alu_result[30]~31_combout ;
wire \M_alu_result[30]~q ;
wire \E_src1[30]~33_combout ;
wire \D_src1_prelim[30]~19_combout ;
wire \E_src1_prelim[30]~q ;
wire \E_src1[30]~34_combout ;
wire \E_src1[30]~35_combout ;
wire \M_shift_rot_result_nxt[30]~19_combout ;
wire \M_shift_rot_result[30]~q ;
wire \W_wr_data[31]~q ;
wire \D_src1_prelim[31]~17_combout ;
wire \E_src1_prelim[31]~q ;
wire \E_src1[31]~31_combout ;
wire \M_shift_rot_result_nxt[31]~17_combout ;
wire \M_shift_rot_result[31]~q ;
wire \av_ld_data_aligned_or_div[31]~q ;
wire \Equal4~14_combout ;
wire \Equal4~15_combout ;
wire \D_ctrl_alu_signed_comparison~0_combout ;
wire \D_ctrl_alu_signed_comparison~1_combout ;
wire \E_ctrl_alu_signed_comparison~q ;
wire \D_src2_imm[31]~0_combout ;
wire \E_src2_imm[31]~q ;
wire \D_src2_prelim[31]~17_combout ;
wire \E_src2_prelim[31]~q ;
wire \E_src2[31]~0_combout ;
wire \Add8~82 ;
wire \Add8~73_sumout ;
wire \E_alu_result[31]~26_combout ;
wire \E_alu_result[31]~27_combout ;
wire \M_alu_result[31]~q ;
wire \M_wr_data_unfiltered[31]~17_combout ;
wire \E_logic_result~0_combout ;
wire \E_logic_result~1_combout ;
wire \E_logic_result~2_combout ;
wire \E_logic_result~3_combout ;
wire \E_logic_result~4_combout ;
wire \E_logic_result~5_combout ;
wire \E_logic_result~6_combout ;
wire \E_logic_result~7_combout ;
wire \E_arith_src2[15]~2_combout ;
wire \E_logic_result~18_combout ;
wire \E_arith_src2[13]~4_combout ;
wire \E_logic_result~14_combout ;
wire \E_arith_src2[11]~6_combout ;
wire \E_logic_result~8_combout ;
wire \E_arith_src2[9]~7_combout ;
wire \E_logic_result~9_combout ;
wire \E_arith_src2[7]~8_combout ;
wire \E_logic_result~10_combout ;
wire \E_arith_src2[5]~0_combout ;
wire \E_logic_result~11_combout ;
wire \E_arith_src2[3]~9_combout ;
wire \D_src1_prelim[3]~13_combout ;
wire \E_src1_prelim[3]~q ;
wire \E_logic_result~12_combout ;
wire \D_src2_prelim[1]~16_combout ;
wire \E_src2_prelim[1]~q ;
wire \E_arith_src2[1]~12_combout ;
wire \E_logic_result~13_combout ;
wire \Add10~130_cout ;
wire \Add10~126_cout ;
wire \Add10~122_cout ;
wire \Add10~118_cout ;
wire \Add10~114_cout ;
wire \Add10~110_cout ;
wire \Add10~106_cout ;
wire \Add10~102_cout ;
wire \Add10~98_cout ;
wire \Add10~94_cout ;
wire \Add10~90_cout ;
wire \Add10~86_cout ;
wire \Add10~82_cout ;
wire \Add10~78_cout ;
wire \Add10~74_cout ;
wire \Add10~70_cout ;
wire \Add10~66_cout ;
wire \Add10~62_cout ;
wire \Add10~58_cout ;
wire \Add10~54_cout ;
wire \Add10~50_cout ;
wire \Add10~46_cout ;
wire \Add10~42_cout ;
wire \Add10~38_cout ;
wire \Add10~34_cout ;
wire \Add10~30_cout ;
wire \Add10~26_cout ;
wire \Add10~22_cout ;
wire \Add10~18_cout ;
wire \Add10~14_cout ;
wire \Add10~10_cout ;
wire \Add10~6_cout ;
wire \Add10~1_sumout ;
wire \Add8~74 ;
wire \Add8~61_sumout ;
wire \D_ctrl_break~1_combout ;
wire \E_ctrl_break~q ;
wire \D_ctrl_exception~1_combout ;
wire \D_ctrl_exception~combout ;
wire \E_ctrl_exception~q ;
wire \D_ctrl_crst~1_combout ;
wire \E_ctrl_crst~q ;
wire \E_iw[6]~q ;
wire \E_iw[7]~q ;
wire \E_iw[8]~q ;
wire \Equal107~2_combout ;
wire \E_ctrl_wrctl_inst~q ;
wire \E_op_eret~1_combout ;
wire \M_status_reg_pie_inst_nxt~0_combout ;
wire \E_wrctl_estatus~combout ;
wire \M_estatus_reg_pie_inst_nxt~0_combout ;
wire \M_estatus_reg_pie~q ;
wire \E_wrctl_bstatus~combout ;
wire \M_bstatus_reg_pie_inst_nxt~0_combout ;
wire \M_bstatus_reg_pie~q ;
wire \M_status_reg_pie_inst_nxt~1_combout ;
wire \M_status_reg_pie_inst_nxt~2_combout ;
wire \M_status_reg_pie_inst_nxt~3_combout ;
wire \M_status_reg_pie~q ;
wire \D_control_reg_rddata_muxed[0]~1_combout ;
wire \E_control_reg_rddata[0]~q ;
wire \Add8~65_sumout ;
wire \E_wrctl_data_bstatus_reg_pie~0_combout ;
wire \E_wrctl_data_bstatus_reg_pie~1_combout ;
wire \E_wrctl_data_bstatus_reg_pie~2_combout ;
wire \M_alu_result[0]~q ;
wire \M_ld_align_sh8~combout ;
wire \av_ld_byte0_data[1]~7_combout ;
wire \av_ld_data_aligned_or_div[1]~q ;
wire \M_wr_data_unfiltered[1]~9_combout ;
wire \E_stb_data[1]~12_combout ;
wire \Add8~69_sumout ;
wire \M_ienable_reg_irq16~1_combout ;
wire \M_ienable_reg_irq16~0_combout ;
wire \M_ienable_reg_irq1~q ;
wire \M_ipending_reg_irq1_nxt~combout ;
wire \M_ipending_reg_irq1~q ;
wire \D_control_reg_rddata_muxed[1]~2_combout ;
wire \E_control_reg_rddata[1]~q ;
wire \E_wrctl_data_ienable_reg_irq1~0_combout ;
wire \E_wrctl_data_ienable_reg_irq1~1_combout ;
wire \M_alu_result[1]~q ;
wire \M_ld_align_sh16~combout ;
wire \av_ld_byte0_data[3]~5_combout ;
wire \av_ld_data_aligned_or_div[3]~q ;
wire \M_wr_data_unfiltered[3]~8_combout ;
wire \E_src1[3]~23_combout ;
wire \M_shift_rot_result_nxt[3]~14_combout ;
wire \M_shift_rot_result[3]~q ;
wire \M_shift_rot_result_nxt[2]~15_combout ;
wire \M_shift_rot_result[2]~q ;
wire \M_shift_rot_result_nxt[1]~16_combout ;
wire \M_shift_rot_result[1]~q ;
wire \M_shift_rot_result_nxt[0]~0_combout ;
wire \M_shift_rot_result[0]~q ;
wire \M_wr_data_unfiltered[0]~10_combout ;
wire \D_src2_prelim[0]~0_combout ;
wire \E_src2_prelim[0]~q ;
wire \E_stb_data[0]~1_combout ;
wire \E_arith_src2[0]~11_combout ;
wire \M_shift_rot_cnt[0]~q ;
wire \M_shift_rot_cnt_nxt[0]~0_combout ;
wire \M_shift_rot_cnt[1]~q ;
wire \M_shift_rot_cnt_nxt[1]~1_combout ;
wire \E_arith_src2[2]~10_combout ;
wire \M_shift_rot_cnt[2]~q ;
wire \M_shift_rot_cnt_nxt[2]~2_combout ;
wire \E_arith_src2[4]~1_combout ;
wire \M_shift_rot_cnt[4]~q ;
wire \Add9~0_combout ;
wire \M_shift_rot_cnt_nxt[3]~4_combout ;
wire \M_shift_rot_cnt[3]~q ;
wire \M_shift_rot_cnt_nxt[4]~3_combout ;
wire \Equal198~0_combout ;
wire \M_shift_rot_stall_nxt~0_combout ;
wire \M_shift_rot_stall~q ;
wire \W_stall~0_combout ;
wire \W_stall~combout ;
wire \D_iw[14]~q ;
wire \E_iw[14]~q ;
wire \E_hbreak_req~combout ;
wire \E_iw[21]~q ;
wire \E_br_mispredict~0_combout ;
wire \E_ctrl_br_cond_nxt~0_combout ;
wire \E_ctrl_br_cond_nxt~1_combout ;
wire \E_ctrl_br_cond~q ;
wire \Equal4~11_combout ;
wire \Equal4~13_combout ;
wire \D_ctrl_flush_pipe_always~1_combout ;
wire \D_ctrl_flush_pipe_always~0_combout ;
wire \E_ctrl_flush_pipe_always~q ;
wire \M_pipe_flush_nxt~0_combout ;
wire \M_pipe_flush~q ;
wire \D_ctrl_br~0_combout ;
wire \Equal4~12_combout ;
wire \D_ctrl_jmp_indirect~0_combout ;
wire \E_ctrl_jmp_indirect~q ;
wire \E_ctrl_jmp_direct~q ;
wire \M_pipe_flush_waddr[7]~0_combout ;
wire \Add3~57_sumout ;
wire \Add0~37_sumout ;
wire \D_br_taken_waddr_partial[0]~q ;
wire \D_pc_plus_one[0]~q ;
wire \D_br_pred_not_taken~combout ;
wire \E_extra_pc[0]~q ;
wire \M_pipe_flush_waddr[7]~1_combout ;
wire \M_pipe_flush_waddr_nxt[0]~0_combout ;
wire \M_pipe_flush_waddr_nxt[0]~1_combout ;
wire \D_pc[0]~q ;
wire \E_pc[0]~q ;
wire \M_pipe_flush_waddr[7]~2_combout ;
wire \M_pipe_flush_waddr[0]~q ;
wire \F_ic_data_rd_addr_nxt[0]~0_combout ;
wire \F_ic_data_rd_addr_nxt[0]~1_combout ;
wire \F_pc[0]~q ;
wire \Add3~58 ;
wire \Add3~53_sumout ;
wire \Add0~38 ;
wire \Add0~33_sumout ;
wire \D_br_taken_waddr_partial[1]~q ;
wire \D_pc_plus_one[1]~q ;
wire \E_extra_pc[1]~q ;
wire \M_pipe_flush_waddr_nxt[1]~2_combout ;
wire \M_pipe_flush_waddr_nxt[1]~3_combout ;
wire \D_pc[1]~q ;
wire \E_pc[1]~q ;
wire \M_pipe_flush_waddr[1]~q ;
wire \F_ic_data_rd_addr_nxt[1]~2_combout ;
wire \F_pc[1]~q ;
wire \Add3~54 ;
wire \Add3~5_sumout ;
wire \Add0~34 ;
wire \Add0~5_sumout ;
wire \D_br_taken_waddr_partial[2]~q ;
wire \D_pc_plus_one[2]~q ;
wire \E_extra_pc[2]~q ;
wire \M_pipe_flush_waddr_nxt[2]~4_combout ;
wire \M_pipe_flush_waddr_nxt[2]~5_combout ;
wire \D_pc[2]~q ;
wire \E_pc[2]~q ;
wire \M_pipe_flush_waddr[2]~q ;
wire \F_ic_data_rd_addr_nxt[2]~3_combout ;
wire \F_pc[2]~q ;
wire \F_ic_valid~4_combout ;
wire \F_ic_valid~0_combout ;
wire \D_pc[13]~q ;
wire \E_pc[13]~q ;
wire \Add3~6 ;
wire \Add3~1_sumout ;
wire \Add0~6 ;
wire \Add0~1_sumout ;
wire \D_br_taken_waddr_partial[3]~q ;
wire \D_pc_plus_one[3]~q ;
wire \E_extra_pc[3]~q ;
wire \M_pipe_flush_waddr_nxt[3]~6_combout ;
wire \E_iw[9]~q ;
wire \M_pipe_flush_waddr_nxt[3]~7_combout ;
wire \D_pc[3]~q ;
wire \E_pc[3]~q ;
wire \M_pipe_flush_waddr[3]~q ;
wire \F_ic_tag_rd_addr_nxt[0]~0_combout ;
wire \F_pc[3]~q ;
wire \Add3~2 ;
wire \Add3~9_sumout ;
wire \Add0~2 ;
wire \Add0~9_sumout ;
wire \D_br_taken_waddr_partial[4]~q ;
wire \D_pc_plus_one[4]~q ;
wire \E_extra_pc[4]~q ;
wire \M_pipe_flush_waddr_nxt[4]~8_combout ;
wire \E_iw[10]~q ;
wire \M_pipe_flush_waddr_nxt[4]~9_combout ;
wire \D_pc[4]~q ;
wire \E_pc[4]~q ;
wire \M_pipe_flush_waddr[4]~q ;
wire \F_ic_tag_rd_addr_nxt[1]~1_combout ;
wire \F_pc[4]~q ;
wire \Add3~10 ;
wire \Add3~49_sumout ;
wire \Add0~10 ;
wire \Add0~29_sumout ;
wire \D_br_taken_waddr_partial[5]~q ;
wire \D_pc_plus_one[5]~q ;
wire \E_extra_pc[5]~q ;
wire \M_pipe_flush_waddr_nxt[5]~10_combout ;
wire \M_pipe_flush_waddr_nxt[5]~11_combout ;
wire \D_pc[5]~q ;
wire \E_pc[5]~q ;
wire \M_pipe_flush_waddr[5]~q ;
wire \F_ic_tag_rd_addr_nxt[2]~2_combout ;
wire \F_pc[5]~q ;
wire \Add3~50 ;
wire \Add3~45_sumout ;
wire \Add0~30 ;
wire \Add0~25_sumout ;
wire \D_br_taken_waddr_partial[6]~q ;
wire \D_pc_plus_one[6]~q ;
wire \E_extra_pc[6]~q ;
wire \M_pipe_flush_waddr_nxt[6]~12_combout ;
wire \M_pipe_flush_waddr_nxt[6]~13_combout ;
wire \D_pc[6]~q ;
wire \E_pc[6]~q ;
wire \M_pipe_flush_waddr[6]~q ;
wire \F_ic_tag_rd_addr_nxt[3]~3_combout ;
wire \F_pc[6]~q ;
wire \Add3~46 ;
wire \Add3~41_sumout ;
wire \Add0~26 ;
wire \Add0~21_sumout ;
wire \D_br_taken_waddr_partial[7]~q ;
wire \D_pc_plus_one[7]~q ;
wire \E_extra_pc[7]~q ;
wire \M_pipe_flush_waddr_nxt[7]~14_combout ;
wire \M_pipe_flush_waddr_nxt[7]~15_combout ;
wire \D_pc[7]~q ;
wire \E_pc[7]~q ;
wire \M_pipe_flush_waddr[7]~q ;
wire \F_ic_tag_rd_addr_nxt[4]~4_combout ;
wire \F_pc[7]~q ;
wire \Add3~42 ;
wire \Add3~37_sumout ;
wire \Add0~22 ;
wire \Add0~17_sumout ;
wire \D_br_taken_waddr_partial[8]~q ;
wire \D_pc_plus_one[8]~q ;
wire \E_extra_pc[8]~q ;
wire \M_pipe_flush_waddr_nxt[8]~16_combout ;
wire \M_pipe_flush_waddr_nxt[8]~17_combout ;
wire \D_pc[8]~q ;
wire \E_pc[8]~q ;
wire \M_pipe_flush_waddr[8]~q ;
wire \F_ic_tag_rd_addr_nxt[5]~5_combout ;
wire \F_pc[8]~q ;
wire \Add3~38 ;
wire \Add3~33_sumout ;
wire \Add0~18 ;
wire \Add0~13_sumout ;
wire \D_br_taken_waddr_partial[9]~q ;
wire \D_pc_plus_one[9]~q ;
wire \E_extra_pc[9]~q ;
wire \M_pipe_flush_waddr[7]~3_combout ;
wire \M_pipe_flush_waddr_nxt[9]~23_combout ;
wire \D_pc[9]~q ;
wire \E_pc[9]~q ;
wire \M_pipe_flush_waddr[9]~q ;
wire \F_pc_nxt[9]~3_combout ;
wire \F_pc[9]~q ;
wire \Add3~34 ;
wire \Add3~29_sumout ;
wire \D_pc_plus_one[10]~q ;
wire \Add0~14 ;
wire \Add0~41_sumout ;
wire \D_br_taken_waddr_partial[10]~q ;
wire \Add1~22_cout ;
wire \Add1~17_sumout ;
wire \E_extra_pc[10]~q ;
wire \M_pipe_flush_waddr_nxt[10]~19_combout ;
wire \M_pipe_flush_waddr_nxt[10]~20_combout ;
wire \D_pc[10]~q ;
wire \E_pc[10]~q ;
wire \M_pipe_flush_waddr[10]~q ;
wire \F_pc_nxt[10]~1_combout ;
wire \F_pc[10]~q ;
wire \Add3~30 ;
wire \Add3~25_sumout ;
wire \D_pc_plus_one[11]~q ;
wire \Add1~18 ;
wire \Add1~13_sumout ;
wire \E_extra_pc[11]~q ;
wire \M_pipe_flush_waddr_nxt[11]~24_combout ;
wire \E_iw[17]~q ;
wire \M_pipe_flush_waddr_nxt[11]~25_combout ;
wire \D_pc[11]~q ;
wire \E_pc[11]~q ;
wire \M_pipe_flush_waddr[11]~q ;
wire \F_pc_nxt[11]~4_combout ;
wire \F_pc[11]~q ;
wire \Add3~26 ;
wire \Add3~21_sumout ;
wire \D_pc_plus_one[12]~q ;
wire \Add1~14 ;
wire \Add1~9_sumout ;
wire \E_extra_pc[12]~q ;
wire \M_pipe_flush_waddr_nxt[12]~26_combout ;
wire \E_iw[18]~q ;
wire \M_pipe_flush_waddr_nxt[12]~27_combout ;
wire \D_pc[12]~q ;
wire \E_pc[12]~q ;
wire \M_pipe_flush_waddr[12]~q ;
wire \F_pc_nxt[12]~5_combout ;
wire \F_pc[12]~q ;
wire \Add3~22 ;
wire \Add3~17_sumout ;
wire \D_pc_plus_one[13]~q ;
wire \Add1~10 ;
wire \Add1~5_sumout ;
wire \E_extra_pc[13]~q ;
wire \E_iw[19]~q ;
wire \M_pipe_flush_waddr_nxt[13]~21_combout ;
wire \M_pipe_flush_waddr_nxt[13]~22_combout ;
wire \M_pipe_flush_waddr[13]~q ;
wire \F_pc_nxt[13]~2_combout ;
wire \F_pc[13]~q ;
wire \Add3~18 ;
wire \Add3~13_sumout ;
wire \D_pc_plus_one[14]~q ;
wire \Add1~6 ;
wire \Add1~1_sumout ;
wire \E_extra_pc[14]~q ;
wire \E_iw[20]~q ;
wire \M_pipe_flush_waddr_nxt[14]~18_combout ;
wire \D_pc[14]~q ;
wire \E_pc[14]~q ;
wire \M_pipe_flush_waddr[14]~q ;
wire \F_pc_nxt[14]~0_combout ;
wire \F_pc[14]~q ;
wire \W_valid~0_combout ;
wire \W_valid~q ;
wire \M_ctrl_crst~q ;
wire \W_ctrl_crst~q ;
wire \F_inst_ram_hit~0_combout ;
wire \F_inst_ram_hit~1_combout ;
wire \F_inst_ram_hit~2_combout ;
wire \F_inst_ram_hit~3_combout ;
wire \D_iw_valid~q ;
wire \D_kill~q ;
wire \D_refetch~0_combout ;
wire \F_kill~0_combout ;
wire \F_kill~1_combout ;
wire \F_issue~combout ;
wire \D_issue~q ;
wire \D_valid~combout ;
wire \E_valid_from_D~q ;
wire \E_valid~0_combout ;
wire \latched_oci_tb_hbreak_req_next~0_combout ;
wire \latched_oci_tb_hbreak_req~q ;
wire \F_iw~1_combout ;
wire \D_iw[0]~q ;
wire \Equal4~2_combout ;
wire \Equal4~3_combout ;
wire \Equal4~4_combout ;
wire \D_ctrl_logic~0_combout ;
wire \D_ctrl_logic~combout ;
wire \E_ctrl_logic~q ;
wire \Add8~13_sumout ;
wire \E_wrctl_data_ienable_reg_irq16~0_combout ;
wire \D_control_reg_rddata_muxed[16]~0_combout ;
wire \E_control_reg_rddata[16]~q ;
wire \E_wrctl_data_ienable_reg_irq16~1_combout ;
wire \E_wrctl_data_ienable_reg_irq16~2_combout ;
wire \M_ienable_reg_irq16~q ;
wire \M_ipending_reg_irq16_nxt~0_combout ;
wire \M_ipending_reg_irq16~q ;
wire \intr_req~0_combout ;
wire \F_iw[24]~0_combout ;
wire \D_iw[24]~q ;
wire \D_dst_regnum[2]~1_combout ;
wire \E_dst_regnum[2]~q ;
wire \D_src2_hazard_E~0_combout ;
wire \D_src2_hazard_E~1_combout ;
wire \D_src2_hazard_E~combout ;
wire \E_src2_hazard_M~q ;
wire \E_stb_data[0]~0_combout ;
wire \E_stb_data[0]~2_combout ;
wire \Equal0~0_combout ;
wire \D_ctrl_st~0_combout ;
wire \E_ctrl_st~q ;
wire \d_write_nxt~combout ;
wire \Add8~1_sumout ;
wire \E_alu_result[5]~1_combout ;
wire \E_alu_result[5]~2_combout ;
wire \Add8~5_sumout ;
wire \E_alu_result[4]~3_combout ;
wire \E_alu_result[4]~4_combout ;
wire \Add8~9_sumout ;
wire \E_alu_result[6]~64_combout ;
wire \E_alu_result[6]~5_combout ;
wire \Add8~17_sumout ;
wire \E_alu_result[15]~6_combout ;
wire \E_alu_result[15]~7_combout ;
wire \Add8~21_sumout ;
wire \E_arith_src2[14]~3_combout ;
wire \E_alu_result[14]~8_combout ;
wire \E_alu_result[14]~9_combout ;
wire \Add8~25_sumout ;
wire \E_alu_result[13]~10_combout ;
wire \E_alu_result[13]~11_combout ;
wire \Add8~29_sumout ;
wire \E_arith_src2[12]~5_combout ;
wire \E_alu_result[12]~12_combout ;
wire \E_alu_result[12]~13_combout ;
wire \Add8~33_sumout ;
wire \E_alu_result[11]~14_combout ;
wire \E_alu_result[11]~15_combout ;
wire \Add8~37_sumout ;
wire \E_alu_result[10]~60_combout ;
wire \E_alu_result[10]~16_combout ;
wire \Add8~41_sumout ;
wire \E_alu_result[9]~17_combout ;
wire \E_alu_result[9]~18_combout ;
wire \Add8~45_sumout ;
wire \E_alu_result[8]~56_combout ;
wire \E_alu_result[8]~19_combout ;
wire \Add8~49_sumout ;
wire \E_alu_result[7]~20_combout ;
wire \E_alu_result[7]~21_combout ;
wire \Add8~53_sumout ;
wire \E_alu_result[3]~22_combout ;
wire \E_alu_result[3]~23_combout ;
wire \Add8~57_sumout ;
wire \E_alu_result[2]~24_combout ;
wire \E_alu_result[2]~25_combout ;
wire \d_read_nxt~combout ;
wire \M_ctrl_break~q ;
wire \M_iw[11]~q ;
wire \M_iw[1]~q ;
wire \M_iw[0]~q ;
wire \M_iw[16]~q ;
wire \M_iw[15]~q ;
wire \M_iw[14]~q ;
wire \M_iw[13]~q ;
wire \M_iw[12]~q ;
wire \hbreak_enabled~0_combout ;
wire \M_iw[5]~q ;
wire \M_iw[2]~q ;
wire \hbreak_enabled~1_combout ;
wire \hbreak_enabled~2_combout ;
wire \hbreak_enabled~3_combout ;
wire \F_ic_fill_same_tag_line~0_combout ;
wire \F_ic_fill_same_tag_line~1_combout ;
wire \F_ic_fill_same_tag_line~2_combout ;
wire \F_ic_fill_same_tag_line~3_combout ;
wire \F_ic_fill_same_tag_line~4_combout ;
wire \F_ic_fill_same_tag_line~5_combout ;
wire \F_ic_fill_same_tag_line~combout ;
wire \D_ic_fill_same_tag_line~q ;
wire \E_ctrl_invalidate_i~0_combout ;
wire \E_ctrl_invalidate_i~1_combout ;
wire \M_ctrl_invalidate_i~q ;
wire \ic_fill_prevent_refill_nxt~combout ;
wire \ic_fill_prevent_refill~q ;
wire \D_ic_fill_starting~0_combout ;
wire \ic_fill_initial_offset[2]~q ;
wire \ic_fill_initial_offset[0]~q ;
wire \D_ic_fill_starting_d1~q ;
wire \ic_fill_dp_offset_nxt[0]~1_combout ;
wire \i_readdatavalid_d1~q ;
wire \ic_fill_dp_offset_en~0_combout ;
wire \ic_fill_dp_offset[0]~q ;
wire \ic_fill_initial_offset[1]~q ;
wire \ic_fill_dp_offset_nxt[1]~2_combout ;
wire \ic_fill_dp_offset[1]~q ;
wire \ic_fill_dp_offset[2]~q ;
wire \ic_fill_dp_offset_nxt[2]~0_combout ;
wire \ic_fill_active_nxt~0_combout ;
wire \ic_fill_active_nxt~1_combout ;
wire \ic_fill_active~q ;
wire \ic_fill_ap_cnt_nxt[0]~3_combout ;
wire \ic_fill_ap_cnt[2]~0_combout ;
wire \ic_fill_ap_cnt[0]~q ;
wire \ic_fill_ap_cnt_nxt[1]~2_combout ;
wire \ic_fill_ap_cnt[1]~q ;
wire \ic_fill_ap_cnt_nxt[2]~1_combout ;
wire \ic_fill_ap_cnt[2]~q ;
wire \ic_fill_ap_cnt_nxt[3]~0_combout ;
wire \ic_fill_ap_cnt[3]~q ;
wire \i_read_nxt~0_combout ;
wire \i_read_nxt~1_combout ;
wire \ic_tag_wraddress_nxt~0_combout ;
wire \ic_tag_wraddress_nxt~1_combout ;
wire \ic_tag_wraddress_nxt~2_combout ;
wire \ic_tag_wraddress_nxt~3_combout ;
wire \ic_tag_wraddress_nxt~4_combout ;
wire \ic_tag_wraddress_nxt~5_combout ;
wire \ic_fill_ap_offset_nxt[0]~0_combout ;
wire \ic_fill_ap_offset_nxt[1]~1_combout ;
wire \ic_fill_ap_offset_nxt[2]~2_combout ;
wire \E_mem_byte_en~0_combout ;
wire \E_mem_byte_en[2]~1_combout ;
wire \E_mem_byte_en[1]~2_combout ;
wire \E_st_data[24]~0_combout ;
wire \E_mem_byte_en[3]~3_combout ;
wire \E_st_data[29]~1_combout ;
wire \E_st_data[28]~2_combout ;
wire \E_st_data[30]~3_combout ;
wire \E_st_data[31]~4_combout ;
wire \E_st_data[31]~5_combout ;
wire \E_st_data[27]~6_combout ;
wire \E_st_data[26]~7_combout ;
wire \E_st_data[25]~8_combout ;


processor_processor_cpu_register_bank_a_module processor_cpu_register_bank_a(
	.q_b_5(\processor_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[5] ),
	.q_b_4(\processor_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[4] ),
	.q_b_6(\processor_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[6] ),
	.q_b_16(\processor_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[16] ),
	.q_b_15(\processor_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[15] ),
	.q_b_14(\processor_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[14] ),
	.q_b_13(\processor_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[13] ),
	.q_b_12(\processor_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[12] ),
	.q_b_11(\processor_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[11] ),
	.q_b_10(\processor_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[10] ),
	.q_b_9(\processor_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[9] ),
	.q_b_8(\processor_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[8] ),
	.q_b_7(\processor_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[7] ),
	.q_b_3(\processor_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[3] ),
	.q_b_2(\processor_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[2] ),
	.q_b_0(\processor_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[0] ),
	.q_b_29(\processor_cpu_ic_data|the_altsyncram|auto_generated|q_b[29] ),
	.q_b_27(\processor_cpu_ic_data|the_altsyncram|auto_generated|q_b[27] ),
	.q_b_28(\processor_cpu_ic_data|the_altsyncram|auto_generated|q_b[28] ),
	.q_b_30(\processor_cpu_ic_data|the_altsyncram|auto_generated|q_b[30] ),
	.q_b_31(\processor_cpu_ic_data|the_altsyncram|auto_generated|q_b[31] ),
	.q_b_1(\processor_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[1] ),
	.q_b_311(\processor_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[31] ),
	.q_b_17(\processor_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[17] ),
	.q_b_301(\processor_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[30] ),
	.q_b_18(\processor_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[18] ),
	.q_b_291(\processor_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[29] ),
	.q_b_19(\processor_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[19] ),
	.q_b_281(\processor_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[28] ),
	.q_b_24(\processor_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[24] ),
	.q_b_21(\processor_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[21] ),
	.q_b_20(\processor_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[20] ),
	.q_b_22(\processor_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[22] ),
	.q_b_23(\processor_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[23] ),
	.q_b_271(\processor_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[27] ),
	.q_b_26(\processor_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[26] ),
	.q_b_25(\processor_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[25] ),
	.W_stall(\W_stall~combout ),
	.M_wr_data_unfiltered_5(\M_wr_data_unfiltered[5]~0_combout ),
	.M_wr_data_unfiltered_15(\M_wr_data_unfiltered[15]~1_combout ),
	.M_wr_data_unfiltered_14(\M_wr_data_unfiltered[14]~2_combout ),
	.M_wr_data_unfiltered_13(\M_wr_data_unfiltered[13]~3_combout ),
	.M_wr_data_unfiltered_12(\M_wr_data_unfiltered[12]~4_combout ),
	.M_wr_data_unfiltered_11(\M_wr_data_unfiltered[11]~5_combout ),
	.M_wr_data_unfiltered_9(\M_wr_data_unfiltered[9]~6_combout ),
	.M_wr_data_unfiltered_7(\M_wr_data_unfiltered[7]~7_combout ),
	.M_wr_data_unfiltered_3(\M_wr_data_unfiltered[3]~8_combout ),
	.M_wr_data_unfiltered_1(\M_wr_data_unfiltered[1]~9_combout ),
	.M_wr_data_unfiltered_0(\M_wr_data_unfiltered[0]~10_combout ),
	.M_dst_regnum_4(\M_dst_regnum[4]~q ),
	.M_wr_dst_reg(\M_wr_dst_reg~q ),
	.M_dst_regnum_0(\M_dst_regnum[0]~q ),
	.M_dst_regnum_1(\M_dst_regnum[1]~q ),
	.M_dst_regnum_2(\M_dst_regnum[2]~q ),
	.M_dst_regnum_3(\M_dst_regnum[3]~q ),
	.M_wr_data_unfiltered_4(\M_wr_data_unfiltered[4]~11_combout ),
	.M_wr_data_unfiltered_6(\M_wr_data_unfiltered[6]~12_combout ),
	.M_wr_data_unfiltered_16(\M_wr_data_unfiltered[16]~13_combout ),
	.M_wr_data_unfiltered_10(\M_wr_data_unfiltered[10]~14_combout ),
	.M_wr_data_unfiltered_8(\M_wr_data_unfiltered[8]~15_combout ),
	.M_wr_data_unfiltered_2(\M_wr_data_unfiltered[2]~16_combout ),
	.M_wr_data_unfiltered_31(\M_wr_data_unfiltered[31]~17_combout ),
	.M_wr_data_unfiltered_17(\M_wr_data_unfiltered[17]~18_combout ),
	.M_wr_data_unfiltered_30(\M_wr_data_unfiltered[30]~19_combout ),
	.M_wr_data_unfiltered_29(\M_wr_data_unfiltered[29]~20_combout ),
	.M_wr_data_unfiltered_21(\M_wr_data_unfiltered[21]~21_combout ),
	.M_wr_data_unfiltered_19(\M_wr_data_unfiltered[19]~22_combout ),
	.M_wr_data_unfiltered_18(\M_wr_data_unfiltered[18]~23_combout ),
	.M_wr_data_unfiltered_23(\M_wr_data_unfiltered[23]~24_combout ),
	.M_wr_data_unfiltered_27(\M_wr_data_unfiltered[27]~25_combout ),
	.M_wr_data_unfiltered_25(\M_wr_data_unfiltered[25]~26_combout ),
	.M_wr_data_unfiltered_24(\M_wr_data_unfiltered[24]~27_combout ),
	.M_wr_data_unfiltered_20(\M_wr_data_unfiltered[20]~28_combout ),
	.M_wr_data_unfiltered_28(\M_wr_data_unfiltered[28]~29_combout ),
	.M_wr_data_unfiltered_22(\M_wr_data_unfiltered[22]~30_combout ),
	.M_wr_data_unfiltered_26(\M_wr_data_unfiltered[26]~31_combout ),
	.clk_clk(clk_clk));

processor_processor_cpu_ic_tag_module processor_cpu_ic_tag(
	.q_b_5(\processor_cpu_ic_tag|the_altsyncram|auto_generated|q_b[5] ),
	.q_b_1(\processor_cpu_ic_tag|the_altsyncram|auto_generated|q_b[1] ),
	.q_b_4(\processor_cpu_ic_tag|the_altsyncram|auto_generated|q_b[4] ),
	.q_b_0(\processor_cpu_ic_tag|the_altsyncram|auto_generated|q_b[0] ),
	.q_b_2(\processor_cpu_ic_tag|the_altsyncram|auto_generated|q_b[2] ),
	.q_b_3(\processor_cpu_ic_tag|the_altsyncram|auto_generated|q_b[3] ),
	.q_b_11(\processor_cpu_ic_tag|the_altsyncram|auto_generated|q_b[11] ),
	.q_b_13(\processor_cpu_ic_tag|the_altsyncram|auto_generated|q_b[13] ),
	.q_b_10(\processor_cpu_ic_tag|the_altsyncram|auto_generated|q_b[10] ),
	.q_b_12(\processor_cpu_ic_tag|the_altsyncram|auto_generated|q_b[12] ),
	.ic_tag_wraddress_0(\ic_tag_wraddress[0]~q ),
	.ic_fill_valid_bits_5(\ic_fill_valid_bits[5]~q ),
	.ic_fill_valid_bits_7(\ic_fill_valid_bits[7]~q ),
	.ic_fill_valid_bits_4(\ic_fill_valid_bits[4]~q ),
	.q_b_7(\processor_cpu_ic_tag|the_altsyncram|auto_generated|q_b[7] ),
	.q_b_9(\processor_cpu_ic_tag|the_altsyncram|auto_generated|q_b[9] ),
	.q_b_6(\processor_cpu_ic_tag|the_altsyncram|auto_generated|q_b[6] ),
	.q_b_8(\processor_cpu_ic_tag|the_altsyncram|auto_generated|q_b[8] ),
	.ic_fill_valid_bits_6(\ic_fill_valid_bits[6]~q ),
	.ic_fill_valid_bits_1(\ic_fill_valid_bits[1]~q ),
	.ic_fill_valid_bits_3(\ic_fill_valid_bits[3]~q ),
	.ic_fill_valid_bits_0(\ic_fill_valid_bits[0]~q ),
	.ic_fill_valid_bits_2(\ic_fill_valid_bits[2]~q ),
	.W_stall(\W_stall~combout ),
	.ic_fill_tag_5(ic_fill_tag_5),
	.ic_fill_tag_4(ic_fill_tag_4),
	.ic_fill_tag_3(ic_fill_tag_3),
	.ic_fill_tag_2(ic_fill_tag_2),
	.ic_fill_tag_1(ic_fill_tag_1),
	.ic_fill_tag_0(ic_fill_tag_0),
	.F_ic_tag_rd_addr_nxt_0(\F_ic_tag_rd_addr_nxt[0]~0_combout ),
	.F_ic_tag_rd_addr_nxt_1(\F_ic_tag_rd_addr_nxt[1]~1_combout ),
	.F_ic_tag_rd_addr_nxt_2(\F_ic_tag_rd_addr_nxt[2]~2_combout ),
	.F_ic_tag_rd_addr_nxt_3(\F_ic_tag_rd_addr_nxt[3]~3_combout ),
	.F_ic_tag_rd_addr_nxt_4(\F_ic_tag_rd_addr_nxt[4]~4_combout ),
	.F_ic_tag_rd_addr_nxt_5(\F_ic_tag_rd_addr_nxt[5]~5_combout ),
	.ic_tag_wren(\ic_tag_wren~combout ),
	.ic_tag_wraddress_1(\ic_tag_wraddress[1]~q ),
	.ic_tag_wraddress_2(\ic_tag_wraddress[2]~q ),
	.ic_tag_wraddress_3(\ic_tag_wraddress[3]~q ),
	.ic_tag_wraddress_4(\ic_tag_wraddress[4]~q ),
	.ic_tag_wraddress_5(\ic_tag_wraddress[5]~q ),
	.clk_clk(clk_clk));

processor_processor_cpu_ic_data_module processor_cpu_ic_data(
	.q_b_24(\processor_cpu_ic_data|the_altsyncram|auto_generated|q_b[24] ),
	.q_b_0(\processor_cpu_ic_data|the_altsyncram|auto_generated|q_b[0] ),
	.q_b_1(\processor_cpu_ic_data|the_altsyncram|auto_generated|q_b[1] ),
	.q_b_2(\processor_cpu_ic_data|the_altsyncram|auto_generated|q_b[2] ),
	.q_b_3(\processor_cpu_ic_data|the_altsyncram|auto_generated|q_b[3] ),
	.q_b_4(\processor_cpu_ic_data|the_altsyncram|auto_generated|q_b[4] ),
	.q_b_5(\processor_cpu_ic_data|the_altsyncram|auto_generated|q_b[5] ),
	.q_b_22(\processor_cpu_ic_data|the_altsyncram|auto_generated|q_b[22] ),
	.q_b_23(\processor_cpu_ic_data|the_altsyncram|auto_generated|q_b[23] ),
	.q_b_25(\processor_cpu_ic_data|the_altsyncram|auto_generated|q_b[25] ),
	.q_b_26(\processor_cpu_ic_data|the_altsyncram|auto_generated|q_b[26] ),
	.q_b_14(\processor_cpu_ic_data|the_altsyncram|auto_generated|q_b[14] ),
	.q_b_12(\processor_cpu_ic_data|the_altsyncram|auto_generated|q_b[12] ),
	.q_b_11(\processor_cpu_ic_data|the_altsyncram|auto_generated|q_b[11] ),
	.q_b_16(\processor_cpu_ic_data|the_altsyncram|auto_generated|q_b[16] ),
	.q_b_15(\processor_cpu_ic_data|the_altsyncram|auto_generated|q_b[15] ),
	.q_b_13(\processor_cpu_ic_data|the_altsyncram|auto_generated|q_b[13] ),
	.q_b_21(\processor_cpu_ic_data|the_altsyncram|auto_generated|q_b[21] ),
	.q_b_29(\processor_cpu_ic_data|the_altsyncram|auto_generated|q_b[29] ),
	.q_b_27(\processor_cpu_ic_data|the_altsyncram|auto_generated|q_b[27] ),
	.q_b_28(\processor_cpu_ic_data|the_altsyncram|auto_generated|q_b[28] ),
	.q_b_30(\processor_cpu_ic_data|the_altsyncram|auto_generated|q_b[30] ),
	.q_b_31(\processor_cpu_ic_data|the_altsyncram|auto_generated|q_b[31] ),
	.q_b_10(\processor_cpu_ic_data|the_altsyncram|auto_generated|q_b[10] ),
	.q_b_6(\processor_cpu_ic_data|the_altsyncram|auto_generated|q_b[6] ),
	.q_b_8(\processor_cpu_ic_data|the_altsyncram|auto_generated|q_b[8] ),
	.q_b_7(\processor_cpu_ic_data|the_altsyncram|auto_generated|q_b[7] ),
	.q_b_20(\processor_cpu_ic_data|the_altsyncram|auto_generated|q_b[20] ),
	.q_b_19(\processor_cpu_ic_data|the_altsyncram|auto_generated|q_b[19] ),
	.q_b_18(\processor_cpu_ic_data|the_altsyncram|auto_generated|q_b[18] ),
	.q_b_17(\processor_cpu_ic_data|the_altsyncram|auto_generated|q_b[17] ),
	.q_b_9(\processor_cpu_ic_data|the_altsyncram|auto_generated|q_b[9] ),
	.W_stall(\W_stall~combout ),
	.ic_fill_line_5(ic_fill_line_5),
	.i_readdatavalid_d1(\i_readdatavalid_d1~q ),
	.i_readdata_d1_24(\i_readdata_d1[24]~q ),
	.ic_fill_dp_offset_0(\ic_fill_dp_offset[0]~q ),
	.ic_fill_dp_offset_1(\ic_fill_dp_offset[1]~q ),
	.ic_fill_dp_offset_2(\ic_fill_dp_offset[2]~q ),
	.ic_fill_line_0(ic_fill_line_0),
	.ic_fill_line_1(ic_fill_line_1),
	.ic_fill_line_2(ic_fill_line_2),
	.ic_fill_line_3(ic_fill_line_3),
	.ic_fill_line_4(ic_fill_line_4),
	.F_ic_data_rd_addr_nxt_0(\F_ic_data_rd_addr_nxt[0]~1_combout ),
	.F_ic_data_rd_addr_nxt_1(\F_ic_data_rd_addr_nxt[1]~2_combout ),
	.F_ic_data_rd_addr_nxt_2(\F_ic_data_rd_addr_nxt[2]~3_combout ),
	.F_ic_tag_rd_addr_nxt_0(\F_ic_tag_rd_addr_nxt[0]~0_combout ),
	.F_ic_tag_rd_addr_nxt_1(\F_ic_tag_rd_addr_nxt[1]~1_combout ),
	.F_ic_tag_rd_addr_nxt_2(\F_ic_tag_rd_addr_nxt[2]~2_combout ),
	.F_ic_tag_rd_addr_nxt_3(\F_ic_tag_rd_addr_nxt[3]~3_combout ),
	.F_ic_tag_rd_addr_nxt_4(\F_ic_tag_rd_addr_nxt[4]~4_combout ),
	.F_ic_tag_rd_addr_nxt_5(\F_ic_tag_rd_addr_nxt[5]~5_combout ),
	.i_readdata_d1_0(\i_readdata_d1[0]~q ),
	.i_readdata_d1_1(\i_readdata_d1[1]~q ),
	.i_readdata_d1_2(\i_readdata_d1[2]~q ),
	.i_readdata_d1_3(\i_readdata_d1[3]~q ),
	.i_readdata_d1_4(\i_readdata_d1[4]~q ),
	.i_readdata_d1_5(\i_readdata_d1[5]~q ),
	.i_readdata_d1_22(\i_readdata_d1[22]~q ),
	.i_readdata_d1_23(\i_readdata_d1[23]~q ),
	.i_readdata_d1_25(\i_readdata_d1[25]~q ),
	.i_readdata_d1_26(\i_readdata_d1[26]~q ),
	.i_readdata_d1_14(\i_readdata_d1[14]~q ),
	.i_readdata_d1_12(\i_readdata_d1[12]~q ),
	.i_readdata_d1_11(\i_readdata_d1[11]~q ),
	.i_readdata_d1_16(\i_readdata_d1[16]~q ),
	.i_readdata_d1_15(\i_readdata_d1[15]~q ),
	.i_readdata_d1_13(\i_readdata_d1[13]~q ),
	.i_readdata_d1_21(\i_readdata_d1[21]~q ),
	.i_readdata_d1_29(\i_readdata_d1[29]~q ),
	.i_readdata_d1_27(\i_readdata_d1[27]~q ),
	.i_readdata_d1_28(\i_readdata_d1[28]~q ),
	.i_readdata_d1_30(\i_readdata_d1[30]~q ),
	.i_readdata_d1_31(\i_readdata_d1[31]~q ),
	.i_readdata_d1_10(\i_readdata_d1[10]~q ),
	.i_readdata_d1_6(\i_readdata_d1[6]~q ),
	.i_readdata_d1_8(\i_readdata_d1[8]~q ),
	.i_readdata_d1_7(\i_readdata_d1[7]~q ),
	.i_readdata_d1_20(\i_readdata_d1[20]~q ),
	.i_readdata_d1_19(\i_readdata_d1[19]~q ),
	.i_readdata_d1_18(\i_readdata_d1[18]~q ),
	.i_readdata_d1_17(\i_readdata_d1[17]~q ),
	.i_readdata_d1_9(\i_readdata_d1[9]~q ),
	.clk_clk(clk_clk));

processor_processor_cpu_nios2_oci the_processor_cpu_nios2_oci(
	.readdata_0(readdata_0),
	.readdata_16(readdata_16),
	.readdata_8(readdata_8),
	.readdata_24(readdata_24),
	.readdata_5(readdata_5),
	.readdata_21(readdata_21),
	.readdata_13(readdata_13),
	.readdata_29(readdata_29),
	.readdata_4(readdata_4),
	.readdata_20(readdata_20),
	.readdata_12(readdata_12),
	.readdata_28(readdata_28),
	.readdata_6(readdata_6),
	.readdata_22(readdata_22),
	.readdata_14(readdata_14),
	.readdata_30(readdata_30),
	.readdata_7(readdata_7),
	.readdata_23(readdata_23),
	.readdata_15(readdata_15),
	.readdata_31(readdata_31),
	.readdata_11(readdata_11),
	.readdata_27(readdata_27),
	.readdata_10(readdata_10),
	.readdata_26(readdata_26),
	.readdata_25(readdata_25),
	.readdata_9(readdata_9),
	.readdata_3(readdata_3),
	.readdata_19(readdata_19),
	.readdata_2(readdata_2),
	.readdata_18(readdata_18),
	.readdata_1(readdata_1),
	.readdata_17(readdata_17),
	.sr_0(sr_0),
	.ir_out_0(ir_out_0),
	.ir_out_1(ir_out_1),
	.r_sync_rst(r_sync_rst),
	.d_write(d_write1),
	.saved_grant_0(saved_grant_0),
	.waitrequest(jtag_debug_module_waitrequest),
	.mem_used_1(mem_used_1),
	.hbreak_enabled(hbreak_enabled1),
	.jtag_break(\the_processor_cpu_nios2_oci|the_processor_cpu_nios2_oci_debug|jtag_break~q ),
	.src2_valid(src2_valid),
	.saved_grant_1(saved_grant_1),
	.src0_valid(src0_valid),
	.rf_source_valid(rf_source_valid),
	.oci_single_step_mode(\the_processor_cpu_nios2_oci|the_processor_cpu_nios2_avalon_reg|oci_single_step_mode~q ),
	.address_nxt({src_data_46,src_data_45,src_data_44,src_data_43,src_data_42,src_data_41,src_data_40,src_data_39,src_data_38}),
	.oci_ienable_16(\the_processor_cpu_nios2_oci|the_processor_cpu_nios2_avalon_reg|oci_ienable[16]~q ),
	.r_early_rst(r_early_rst),
	.oci_ienable_1(\the_processor_cpu_nios2_oci|the_processor_cpu_nios2_avalon_reg|oci_ienable[1]~q ),
	.writedata_nxt({src_payload24,src_payload20,src_payload13,src_payload16,src_payload26,src_payload28,src_payload29,src_payload7,src_payload22,src_payload18,src_payload11,src_payload8,src_payload9,src_payload31,src_payload32,src_payload3,src_payload23,src_payload19,src_payload12,src_payload15,
src_payload25,src_payload27,src_payload30,src_payload6,src_payload21,src_payload17,src_payload10,src_payload14,src_payload,src_payload5,src_payload4,src_payload2}),
	.debugaccess_nxt(src_payload1),
	.byteenable_nxt({src_data_35,src_data_34,src_data_33,src_data_32}),
	.altera_internal_jtag(altera_internal_jtag),
	.altera_internal_jtag1(altera_internal_jtag1),
	.state_1(state_1),
	.state_4(state_4),
	.virtual_ir_scan_reg(virtual_ir_scan_reg),
	.state_3(state_3),
	.state_8(state_8),
	.splitter_nodes_receive_1_3(splitter_nodes_receive_1_3),
	.irf_reg_0_2(irf_reg_0_2),
	.irf_reg_1_2(irf_reg_1_2),
	.clk_clk(clk_clk));

processor_processor_cpu_register_bank_b_module processor_cpu_register_bank_b(
	.q_b_0(\processor_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[0] ),
	.q_b_5(\processor_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[5] ),
	.q_b_4(\processor_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[4] ),
	.q_b_6(\processor_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[6] ),
	.q_b_16(\processor_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[16] ),
	.q_b_15(\processor_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[15] ),
	.q_b_14(\processor_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[14] ),
	.q_b_13(\processor_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[13] ),
	.q_b_12(\processor_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[12] ),
	.q_b_11(\processor_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[11] ),
	.q_b_10(\processor_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[10] ),
	.q_b_9(\processor_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[9] ),
	.q_b_8(\processor_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[8] ),
	.q_b_7(\processor_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[7] ),
	.q_b_3(\processor_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[3] ),
	.q_b_2(\processor_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[2] ),
	.q_b_1(\processor_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[1] ),
	.q_b_24(\processor_cpu_ic_data|the_altsyncram|auto_generated|q_b[24] ),
	.q_b_22(\processor_cpu_ic_data|the_altsyncram|auto_generated|q_b[22] ),
	.q_b_23(\processor_cpu_ic_data|the_altsyncram|auto_generated|q_b[23] ),
	.q_b_25(\processor_cpu_ic_data|the_altsyncram|auto_generated|q_b[25] ),
	.q_b_26(\processor_cpu_ic_data|the_altsyncram|auto_generated|q_b[26] ),
	.q_b_31(\processor_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[31] ),
	.q_b_17(\processor_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[17] ),
	.q_b_30(\processor_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[30] ),
	.q_b_241(\processor_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[24] ),
	.q_b_21(\processor_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[21] ),
	.q_b_29(\processor_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[29] ),
	.q_b_20(\processor_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[20] ),
	.q_b_28(\processor_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[28] ),
	.q_b_221(\processor_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[22] ),
	.q_b_18(\processor_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[18] ),
	.q_b_231(\processor_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[23] ),
	.q_b_27(\processor_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[27] ),
	.q_b_261(\processor_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[26] ),
	.q_b_251(\processor_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[25] ),
	.q_b_19(\processor_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[19] ),
	.W_stall(\W_stall~combout ),
	.M_wr_data_unfiltered_5(\M_wr_data_unfiltered[5]~0_combout ),
	.M_wr_data_unfiltered_15(\M_wr_data_unfiltered[15]~1_combout ),
	.M_wr_data_unfiltered_14(\M_wr_data_unfiltered[14]~2_combout ),
	.M_wr_data_unfiltered_13(\M_wr_data_unfiltered[13]~3_combout ),
	.M_wr_data_unfiltered_12(\M_wr_data_unfiltered[12]~4_combout ),
	.M_wr_data_unfiltered_11(\M_wr_data_unfiltered[11]~5_combout ),
	.M_wr_data_unfiltered_9(\M_wr_data_unfiltered[9]~6_combout ),
	.M_wr_data_unfiltered_7(\M_wr_data_unfiltered[7]~7_combout ),
	.M_wr_data_unfiltered_3(\M_wr_data_unfiltered[3]~8_combout ),
	.M_wr_data_unfiltered_1(\M_wr_data_unfiltered[1]~9_combout ),
	.M_wr_data_unfiltered_0(\M_wr_data_unfiltered[0]~10_combout ),
	.M_dst_regnum_4(\M_dst_regnum[4]~q ),
	.M_wr_dst_reg(\M_wr_dst_reg~q ),
	.M_dst_regnum_0(\M_dst_regnum[0]~q ),
	.M_dst_regnum_1(\M_dst_regnum[1]~q ),
	.M_dst_regnum_2(\M_dst_regnum[2]~q ),
	.M_dst_regnum_3(\M_dst_regnum[3]~q ),
	.M_wr_data_unfiltered_4(\M_wr_data_unfiltered[4]~11_combout ),
	.M_wr_data_unfiltered_6(\M_wr_data_unfiltered[6]~12_combout ),
	.M_wr_data_unfiltered_16(\M_wr_data_unfiltered[16]~13_combout ),
	.M_wr_data_unfiltered_10(\M_wr_data_unfiltered[10]~14_combout ),
	.M_wr_data_unfiltered_8(\M_wr_data_unfiltered[8]~15_combout ),
	.M_wr_data_unfiltered_2(\M_wr_data_unfiltered[2]~16_combout ),
	.M_wr_data_unfiltered_31(\M_wr_data_unfiltered[31]~17_combout ),
	.M_wr_data_unfiltered_17(\M_wr_data_unfiltered[17]~18_combout ),
	.M_wr_data_unfiltered_30(\M_wr_data_unfiltered[30]~19_combout ),
	.M_wr_data_unfiltered_29(\M_wr_data_unfiltered[29]~20_combout ),
	.M_wr_data_unfiltered_21(\M_wr_data_unfiltered[21]~21_combout ),
	.M_wr_data_unfiltered_19(\M_wr_data_unfiltered[19]~22_combout ),
	.M_wr_data_unfiltered_18(\M_wr_data_unfiltered[18]~23_combout ),
	.M_wr_data_unfiltered_23(\M_wr_data_unfiltered[23]~24_combout ),
	.M_wr_data_unfiltered_27(\M_wr_data_unfiltered[27]~25_combout ),
	.M_wr_data_unfiltered_25(\M_wr_data_unfiltered[25]~26_combout ),
	.M_wr_data_unfiltered_24(\M_wr_data_unfiltered[24]~27_combout ),
	.M_wr_data_unfiltered_20(\M_wr_data_unfiltered[20]~28_combout ),
	.M_wr_data_unfiltered_28(\M_wr_data_unfiltered[28]~29_combout ),
	.M_wr_data_unfiltered_22(\M_wr_data_unfiltered[22]~30_combout ),
	.M_wr_data_unfiltered_26(\M_wr_data_unfiltered[26]~31_combout ),
	.clk_clk(clk_clk));

dffeas \ic_tag_wraddress[0] (
	.clk(clk_clk),
	.d(\ic_tag_wraddress_nxt~6_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(!clr_break_line1),
	.ena(vcc),
	.q(\ic_tag_wraddress[0]~q ),
	.prn(vcc));
defparam \ic_tag_wraddress[0] .is_wysiwyg = "true";
defparam \ic_tag_wraddress[0] .power_up = "low";

dffeas \ic_fill_valid_bits[5] (
	.clk(clk_clk),
	.d(\ic_fill_valid_bits_nxt~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\ic_tag_clr_valid_bits_nxt~combout ),
	.sload(gnd),
	.ena(\ic_fill_valid_bits_en~combout ),
	.q(\ic_fill_valid_bits[5]~q ),
	.prn(vcc));
defparam \ic_fill_valid_bits[5] .is_wysiwyg = "true";
defparam \ic_fill_valid_bits[5] .power_up = "low";

dffeas \ic_fill_valid_bits[7] (
	.clk(clk_clk),
	.d(\ic_fill_valid_bits_nxt~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\ic_tag_clr_valid_bits_nxt~combout ),
	.sload(gnd),
	.ena(\ic_fill_valid_bits_en~combout ),
	.q(\ic_fill_valid_bits[7]~q ),
	.prn(vcc));
defparam \ic_fill_valid_bits[7] .is_wysiwyg = "true";
defparam \ic_fill_valid_bits[7] .power_up = "low";

dffeas \ic_fill_valid_bits[4] (
	.clk(clk_clk),
	.d(\ic_fill_valid_bits_nxt~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\ic_tag_clr_valid_bits_nxt~combout ),
	.sload(gnd),
	.ena(\ic_fill_valid_bits_en~combout ),
	.q(\ic_fill_valid_bits[4]~q ),
	.prn(vcc));
defparam \ic_fill_valid_bits[4] .is_wysiwyg = "true";
defparam \ic_fill_valid_bits[4] .power_up = "low";

dffeas \ic_fill_valid_bits[6] (
	.clk(clk_clk),
	.d(\ic_fill_valid_bits_nxt~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\ic_tag_clr_valid_bits_nxt~combout ),
	.sload(gnd),
	.ena(\ic_fill_valid_bits_en~combout ),
	.q(\ic_fill_valid_bits[6]~q ),
	.prn(vcc));
defparam \ic_fill_valid_bits[6] .is_wysiwyg = "true";
defparam \ic_fill_valid_bits[6] .power_up = "low";

dffeas \ic_fill_valid_bits[1] (
	.clk(clk_clk),
	.d(\ic_fill_valid_bits_nxt~4_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\ic_tag_clr_valid_bits_nxt~combout ),
	.sload(gnd),
	.ena(\ic_fill_valid_bits_en~combout ),
	.q(\ic_fill_valid_bits[1]~q ),
	.prn(vcc));
defparam \ic_fill_valid_bits[1] .is_wysiwyg = "true";
defparam \ic_fill_valid_bits[1] .power_up = "low";

dffeas \ic_fill_valid_bits[3] (
	.clk(clk_clk),
	.d(\ic_fill_valid_bits_nxt~5_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\ic_tag_clr_valid_bits_nxt~combout ),
	.sload(gnd),
	.ena(\ic_fill_valid_bits_en~combout ),
	.q(\ic_fill_valid_bits[3]~q ),
	.prn(vcc));
defparam \ic_fill_valid_bits[3] .is_wysiwyg = "true";
defparam \ic_fill_valid_bits[3] .power_up = "low";

dffeas \ic_fill_valid_bits[0] (
	.clk(clk_clk),
	.d(\ic_fill_valid_bits_nxt~6_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\ic_tag_clr_valid_bits_nxt~combout ),
	.sload(gnd),
	.ena(\ic_fill_valid_bits_en~combout ),
	.q(\ic_fill_valid_bits[0]~q ),
	.prn(vcc));
defparam \ic_fill_valid_bits[0] .is_wysiwyg = "true";
defparam \ic_fill_valid_bits[0] .power_up = "low";

dffeas \ic_fill_valid_bits[2] (
	.clk(clk_clk),
	.d(\ic_fill_valid_bits_nxt~7_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\ic_tag_clr_valid_bits_nxt~combout ),
	.sload(gnd),
	.ena(\ic_fill_valid_bits_en~combout ),
	.q(\ic_fill_valid_bits[2]~q ),
	.prn(vcc));
defparam \ic_fill_valid_bits[2] .is_wysiwyg = "true";
defparam \ic_fill_valid_bits[2] .power_up = "low";

dffeas \i_readdata_d1[24] (
	.clk(clk_clk),
	.d(i_readdata[24]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_readdata_d1[24]~q ),
	.prn(vcc));
defparam \i_readdata_d1[24] .is_wysiwyg = "true";
defparam \i_readdata_d1[24] .power_up = "low";

dffeas \i_readdata_d1[0] (
	.clk(clk_clk),
	.d(i_readdata[0]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_readdata_d1[0]~q ),
	.prn(vcc));
defparam \i_readdata_d1[0] .is_wysiwyg = "true";
defparam \i_readdata_d1[0] .power_up = "low";

dffeas \i_readdata_d1[1] (
	.clk(clk_clk),
	.d(i_readdata[1]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_readdata_d1[1]~q ),
	.prn(vcc));
defparam \i_readdata_d1[1] .is_wysiwyg = "true";
defparam \i_readdata_d1[1] .power_up = "low";

dffeas \i_readdata_d1[2] (
	.clk(clk_clk),
	.d(i_readdata[2]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_readdata_d1[2]~q ),
	.prn(vcc));
defparam \i_readdata_d1[2] .is_wysiwyg = "true";
defparam \i_readdata_d1[2] .power_up = "low";

dffeas \i_readdata_d1[3] (
	.clk(clk_clk),
	.d(i_readdata[3]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_readdata_d1[3]~q ),
	.prn(vcc));
defparam \i_readdata_d1[3] .is_wysiwyg = "true";
defparam \i_readdata_d1[3] .power_up = "low";

dffeas \i_readdata_d1[4] (
	.clk(clk_clk),
	.d(i_readdata[4]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_readdata_d1[4]~q ),
	.prn(vcc));
defparam \i_readdata_d1[4] .is_wysiwyg = "true";
defparam \i_readdata_d1[4] .power_up = "low";

dffeas \i_readdata_d1[5] (
	.clk(clk_clk),
	.d(i_readdata[5]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_readdata_d1[5]~q ),
	.prn(vcc));
defparam \i_readdata_d1[5] .is_wysiwyg = "true";
defparam \i_readdata_d1[5] .power_up = "low";

dffeas \i_readdata_d1[22] (
	.clk(clk_clk),
	.d(i_readdata[22]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_readdata_d1[22]~q ),
	.prn(vcc));
defparam \i_readdata_d1[22] .is_wysiwyg = "true";
defparam \i_readdata_d1[22] .power_up = "low";

dffeas \i_readdata_d1[23] (
	.clk(clk_clk),
	.d(i_readdata[23]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_readdata_d1[23]~q ),
	.prn(vcc));
defparam \i_readdata_d1[23] .is_wysiwyg = "true";
defparam \i_readdata_d1[23] .power_up = "low";

dffeas \i_readdata_d1[25] (
	.clk(clk_clk),
	.d(i_readdata[25]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_readdata_d1[25]~q ),
	.prn(vcc));
defparam \i_readdata_d1[25] .is_wysiwyg = "true";
defparam \i_readdata_d1[25] .power_up = "low";

dffeas \i_readdata_d1[26] (
	.clk(clk_clk),
	.d(i_readdata[26]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_readdata_d1[26]~q ),
	.prn(vcc));
defparam \i_readdata_d1[26] .is_wysiwyg = "true";
defparam \i_readdata_d1[26] .power_up = "low";

dffeas \i_readdata_d1[14] (
	.clk(clk_clk),
	.d(i_readdata[14]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_readdata_d1[14]~q ),
	.prn(vcc));
defparam \i_readdata_d1[14] .is_wysiwyg = "true";
defparam \i_readdata_d1[14] .power_up = "low";

dffeas ic_tag_clr_valid_bits(
	.clk(clk_clk),
	.d(\ic_tag_clr_valid_bits~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ic_tag_clr_valid_bits~q ),
	.prn(vcc));
defparam ic_tag_clr_valid_bits.is_wysiwyg = "true";
defparam ic_tag_clr_valid_bits.power_up = "low";

cyclonev_lcell_comb ic_tag_wren(
	.dataa(!\i_readdatavalid_d1~q ),
	.datab(!\ic_tag_clr_valid_bits~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_tag_wren~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam ic_tag_wren.extended_lut = "off";
defparam ic_tag_wren.lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam ic_tag_wren.shared_arith = "off";

dffeas \ic_tag_wraddress[1] (
	.clk(clk_clk),
	.d(\ic_tag_wraddress_nxt[1]~8_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ic_tag_wraddress[1]~q ),
	.prn(vcc));
defparam \ic_tag_wraddress[1] .is_wysiwyg = "true";
defparam \ic_tag_wraddress[1] .power_up = "low";

dffeas \ic_tag_wraddress[2] (
	.clk(clk_clk),
	.d(\ic_tag_wraddress_nxt[2]~9_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ic_tag_wraddress[2]~q ),
	.prn(vcc));
defparam \ic_tag_wraddress[2] .is_wysiwyg = "true";
defparam \ic_tag_wraddress[2] .power_up = "low";

dffeas \ic_tag_wraddress[3] (
	.clk(clk_clk),
	.d(\ic_tag_wraddress_nxt[3]~10_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ic_tag_wraddress[3]~q ),
	.prn(vcc));
defparam \ic_tag_wraddress[3] .is_wysiwyg = "true";
defparam \ic_tag_wraddress[3] .power_up = "low";

dffeas \ic_tag_wraddress[4] (
	.clk(clk_clk),
	.d(\ic_tag_wraddress_nxt[4]~11_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ic_tag_wraddress[4]~q ),
	.prn(vcc));
defparam \ic_tag_wraddress[4] .is_wysiwyg = "true";
defparam \ic_tag_wraddress[4] .power_up = "low";

dffeas \ic_tag_wraddress[5] (
	.clk(clk_clk),
	.d(\ic_tag_wraddress_nxt[5]~12_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ic_tag_wraddress[5]~q ),
	.prn(vcc));
defparam \ic_tag_wraddress[5] .is_wysiwyg = "true";
defparam \ic_tag_wraddress[5] .power_up = "low";

dffeas \i_readdata_d1[12] (
	.clk(clk_clk),
	.d(i_readdata[12]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_readdata_d1[12]~q ),
	.prn(vcc));
defparam \i_readdata_d1[12] .is_wysiwyg = "true";
defparam \i_readdata_d1[12] .power_up = "low";

dffeas \i_readdata_d1[11] (
	.clk(clk_clk),
	.d(i_readdata[11]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_readdata_d1[11]~q ),
	.prn(vcc));
defparam \i_readdata_d1[11] .is_wysiwyg = "true";
defparam \i_readdata_d1[11] .power_up = "low";

dffeas \i_readdata_d1[16] (
	.clk(clk_clk),
	.d(i_readdata[16]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_readdata_d1[16]~q ),
	.prn(vcc));
defparam \i_readdata_d1[16] .is_wysiwyg = "true";
defparam \i_readdata_d1[16] .power_up = "low";

dffeas \i_readdata_d1[15] (
	.clk(clk_clk),
	.d(i_readdata[15]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_readdata_d1[15]~q ),
	.prn(vcc));
defparam \i_readdata_d1[15] .is_wysiwyg = "true";
defparam \i_readdata_d1[15] .power_up = "low";

dffeas \i_readdata_d1[13] (
	.clk(clk_clk),
	.d(i_readdata[13]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_readdata_d1[13]~q ),
	.prn(vcc));
defparam \i_readdata_d1[13] .is_wysiwyg = "true";
defparam \i_readdata_d1[13] .power_up = "low";

dffeas \i_readdata_d1[21] (
	.clk(clk_clk),
	.d(i_readdata[21]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_readdata_d1[21]~q ),
	.prn(vcc));
defparam \i_readdata_d1[21] .is_wysiwyg = "true";
defparam \i_readdata_d1[21] .power_up = "low";

dffeas \i_readdata_d1[29] (
	.clk(clk_clk),
	.d(i_readdata[29]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_readdata_d1[29]~q ),
	.prn(vcc));
defparam \i_readdata_d1[29] .is_wysiwyg = "true";
defparam \i_readdata_d1[29] .power_up = "low";

dffeas \i_readdata_d1[27] (
	.clk(clk_clk),
	.d(i_readdata[27]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_readdata_d1[27]~q ),
	.prn(vcc));
defparam \i_readdata_d1[27] .is_wysiwyg = "true";
defparam \i_readdata_d1[27] .power_up = "low";

dffeas \i_readdata_d1[28] (
	.clk(clk_clk),
	.d(i_readdata[28]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_readdata_d1[28]~q ),
	.prn(vcc));
defparam \i_readdata_d1[28] .is_wysiwyg = "true";
defparam \i_readdata_d1[28] .power_up = "low";

dffeas \i_readdata_d1[30] (
	.clk(clk_clk),
	.d(i_readdata[30]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_readdata_d1[30]~q ),
	.prn(vcc));
defparam \i_readdata_d1[30] .is_wysiwyg = "true";
defparam \i_readdata_d1[30] .power_up = "low";

dffeas \i_readdata_d1[31] (
	.clk(clk_clk),
	.d(i_readdata[31]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_readdata_d1[31]~q ),
	.prn(vcc));
defparam \i_readdata_d1[31] .is_wysiwyg = "true";
defparam \i_readdata_d1[31] .power_up = "low";

dffeas \i_readdata_d1[10] (
	.clk(clk_clk),
	.d(i_readdata[10]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_readdata_d1[10]~q ),
	.prn(vcc));
defparam \i_readdata_d1[10] .is_wysiwyg = "true";
defparam \i_readdata_d1[10] .power_up = "low";

dffeas \i_readdata_d1[6] (
	.clk(clk_clk),
	.d(i_readdata[6]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_readdata_d1[6]~q ),
	.prn(vcc));
defparam \i_readdata_d1[6] .is_wysiwyg = "true";
defparam \i_readdata_d1[6] .power_up = "low";

dffeas \i_readdata_d1[8] (
	.clk(clk_clk),
	.d(i_readdata[8]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_readdata_d1[8]~q ),
	.prn(vcc));
defparam \i_readdata_d1[8] .is_wysiwyg = "true";
defparam \i_readdata_d1[8] .power_up = "low";

dffeas \i_readdata_d1[7] (
	.clk(clk_clk),
	.d(i_readdata[7]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_readdata_d1[7]~q ),
	.prn(vcc));
defparam \i_readdata_d1[7] .is_wysiwyg = "true";
defparam \i_readdata_d1[7] .power_up = "low";

dffeas \i_readdata_d1[20] (
	.clk(clk_clk),
	.d(i_readdata[20]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_readdata_d1[20]~q ),
	.prn(vcc));
defparam \i_readdata_d1[20] .is_wysiwyg = "true";
defparam \i_readdata_d1[20] .power_up = "low";

dffeas \i_readdata_d1[19] (
	.clk(clk_clk),
	.d(i_readdata[19]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_readdata_d1[19]~q ),
	.prn(vcc));
defparam \i_readdata_d1[19] .is_wysiwyg = "true";
defparam \i_readdata_d1[19] .power_up = "low";

dffeas \i_readdata_d1[18] (
	.clk(clk_clk),
	.d(i_readdata[18]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_readdata_d1[18]~q ),
	.prn(vcc));
defparam \i_readdata_d1[18] .is_wysiwyg = "true";
defparam \i_readdata_d1[18] .power_up = "low";

dffeas \i_readdata_d1[17] (
	.clk(clk_clk),
	.d(i_readdata[17]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_readdata_d1[17]~q ),
	.prn(vcc));
defparam \i_readdata_d1[17] .is_wysiwyg = "true";
defparam \i_readdata_d1[17] .power_up = "low";

dffeas \i_readdata_d1[9] (
	.clk(clk_clk),
	.d(i_readdata[9]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_readdata_d1[9]~q ),
	.prn(vcc));
defparam \i_readdata_d1[9] .is_wysiwyg = "true";
defparam \i_readdata_d1[9] .power_up = "low";

cyclonev_lcell_comb ic_tag_clr_valid_bits_nxt(
	.dataa(!clr_break_line1),
	.datab(!\M_valid_from_E~q ),
	.datac(!\D_ic_fill_starting~0_combout ),
	.datad(!\M_ctrl_invalidate_i~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_tag_clr_valid_bits_nxt~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam ic_tag_clr_valid_bits_nxt.extended_lut = "off";
defparam ic_tag_clr_valid_bits_nxt.lut_mask = 64'hBFFFBFFFBFFFBFFF;
defparam ic_tag_clr_valid_bits_nxt.shared_arith = "off";

cyclonev_lcell_comb \ic_tag_wraddress_nxt~6 (
	.dataa(!M_alu_result_5),
	.datab(!\M_valid_from_E~q ),
	.datac(!\M_ctrl_invalidate_i~q ),
	.datad(!\M_ctrl_crst~q ),
	.datae(!\ic_tag_wraddress_nxt~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_tag_wraddress_nxt~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_tag_wraddress_nxt~6 .extended_lut = "off";
defparam \ic_tag_wraddress_nxt~6 .lut_mask = 64'hFF7DFFFFFF7DFFFF;
defparam \ic_tag_wraddress_nxt~6 .shared_arith = "off";

cyclonev_lcell_comb \ic_tag_wraddress_nxt[1]~7 (
	.dataa(!clr_break_line1),
	.datab(!\M_valid_from_E~q ),
	.datac(!\M_ctrl_crst~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_tag_wraddress_nxt[1]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_tag_wraddress_nxt[1]~7 .extended_lut = "off";
defparam \ic_tag_wraddress_nxt[1]~7 .lut_mask = 64'hFDFDFDFDFDFDFDFD;
defparam \ic_tag_wraddress_nxt[1]~7 .shared_arith = "off";

cyclonev_lcell_comb \ic_tag_wraddress_nxt[1]~8 (
	.dataa(!M_alu_result_6),
	.datab(!\M_valid_from_E~q ),
	.datac(!\M_ctrl_invalidate_i~q ),
	.datad(!\ic_tag_wraddress_nxt~2_combout ),
	.datae(!\ic_tag_wraddress_nxt[1]~7_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_tag_wraddress_nxt[1]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_tag_wraddress_nxt[1]~8 .extended_lut = "off";
defparam \ic_tag_wraddress_nxt[1]~8 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \ic_tag_wraddress_nxt[1]~8 .shared_arith = "off";

cyclonev_lcell_comb \ic_tag_wraddress_nxt[2]~9 (
	.dataa(!M_alu_result_7),
	.datab(!\M_valid_from_E~q ),
	.datac(!\M_ctrl_invalidate_i~q ),
	.datad(!\ic_tag_wraddress_nxt~3_combout ),
	.datae(!\ic_tag_wraddress_nxt[1]~7_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_tag_wraddress_nxt[2]~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_tag_wraddress_nxt[2]~9 .extended_lut = "off";
defparam \ic_tag_wraddress_nxt[2]~9 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \ic_tag_wraddress_nxt[2]~9 .shared_arith = "off";

cyclonev_lcell_comb \ic_tag_wraddress_nxt[3]~10 (
	.dataa(!M_alu_result_8),
	.datab(!\M_valid_from_E~q ),
	.datac(!\M_ctrl_invalidate_i~q ),
	.datad(!\ic_tag_wraddress_nxt~4_combout ),
	.datae(!\ic_tag_wraddress_nxt[1]~7_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_tag_wraddress_nxt[3]~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_tag_wraddress_nxt[3]~10 .extended_lut = "off";
defparam \ic_tag_wraddress_nxt[3]~10 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \ic_tag_wraddress_nxt[3]~10 .shared_arith = "off";

cyclonev_lcell_comb \ic_tag_wraddress_nxt[4]~11 (
	.dataa(!M_alu_result_9),
	.datab(!\M_valid_from_E~q ),
	.datac(!\M_ctrl_invalidate_i~q ),
	.datad(!\ic_tag_wraddress_nxt~5_combout ),
	.datae(!\ic_tag_wraddress_nxt[1]~7_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_tag_wraddress_nxt[4]~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_tag_wraddress_nxt[4]~11 .extended_lut = "off";
defparam \ic_tag_wraddress_nxt[4]~11 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \ic_tag_wraddress_nxt[4]~11 .shared_arith = "off";

cyclonev_lcell_comb \ic_tag_wraddress_nxt[5]~12 (
	.dataa(!M_alu_result_10),
	.datab(!\M_valid_from_E~q ),
	.datac(!\M_ctrl_invalidate_i~q ),
	.datad(!\ic_tag_wraddress_nxt~0_combout ),
	.datae(!\ic_tag_wraddress_nxt[1]~7_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_tag_wraddress_nxt[5]~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_tag_wraddress_nxt[5]~12 .extended_lut = "off";
defparam \ic_tag_wraddress_nxt[5]~12 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \ic_tag_wraddress_nxt[5]~12 .shared_arith = "off";

cyclonev_lcell_comb \ic_fill_valid_bits_nxt~0 (
	.dataa(!\D_ic_fill_starting_d1~q ),
	.datab(!\ic_fill_dp_offset_nxt[0]~1_combout ),
	.datac(!\ic_fill_dp_offset_nxt[1]~2_combout ),
	.datad(!\ic_fill_dp_offset_nxt[2]~0_combout ),
	.datae(!\ic_fill_valid_bits[5]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_fill_valid_bits_nxt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_fill_valid_bits_nxt~0 .extended_lut = "off";
defparam \ic_fill_valid_bits_nxt~0 .lut_mask = 64'hFBFFFFFFFBFFFFFF;
defparam \ic_fill_valid_bits_nxt~0 .shared_arith = "off";

cyclonev_lcell_comb ic_fill_valid_bits_en(
	.dataa(!\ic_fill_dp_offset_en~0_combout ),
	.datab(!\ic_tag_clr_valid_bits_nxt~combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_fill_valid_bits_en~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam ic_fill_valid_bits_en.extended_lut = "off";
defparam ic_fill_valid_bits_en.lut_mask = 64'h7777777777777777;
defparam ic_fill_valid_bits_en.shared_arith = "off";

cyclonev_lcell_comb \ic_fill_valid_bits_nxt~1 (
	.dataa(!\D_ic_fill_starting_d1~q ),
	.datab(!\ic_fill_dp_offset_nxt[0]~1_combout ),
	.datac(!\ic_fill_dp_offset_nxt[1]~2_combout ),
	.datad(!\ic_fill_dp_offset_nxt[2]~0_combout ),
	.datae(!\ic_fill_valid_bits[7]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_fill_valid_bits_nxt~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_fill_valid_bits_nxt~1 .extended_lut = "off";
defparam \ic_fill_valid_bits_nxt~1 .lut_mask = 64'hBFFFFFFFBFFFFFFF;
defparam \ic_fill_valid_bits_nxt~1 .shared_arith = "off";

cyclonev_lcell_comb \ic_fill_valid_bits_nxt~2 (
	.dataa(!\D_ic_fill_starting_d1~q ),
	.datab(!\ic_fill_dp_offset_nxt[0]~1_combout ),
	.datac(!\ic_fill_dp_offset_nxt[1]~2_combout ),
	.datad(!\ic_fill_dp_offset_nxt[2]~0_combout ),
	.datae(!\ic_fill_valid_bits[4]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_fill_valid_bits_nxt~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_fill_valid_bits_nxt~2 .extended_lut = "off";
defparam \ic_fill_valid_bits_nxt~2 .lut_mask = 64'hFEFFFFFFFEFFFFFF;
defparam \ic_fill_valid_bits_nxt~2 .shared_arith = "off";

cyclonev_lcell_comb \ic_fill_valid_bits_nxt~3 (
	.dataa(!\D_ic_fill_starting_d1~q ),
	.datab(!\ic_fill_dp_offset_nxt[0]~1_combout ),
	.datac(!\ic_fill_dp_offset_nxt[1]~2_combout ),
	.datad(!\ic_fill_dp_offset_nxt[2]~0_combout ),
	.datae(!\ic_fill_valid_bits[6]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_fill_valid_bits_nxt~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_fill_valid_bits_nxt~3 .extended_lut = "off";
defparam \ic_fill_valid_bits_nxt~3 .lut_mask = 64'hEFFFFFFFEFFFFFFF;
defparam \ic_fill_valid_bits_nxt~3 .shared_arith = "off";

cyclonev_lcell_comb \ic_fill_valid_bits_nxt~4 (
	.dataa(!\D_ic_fill_starting_d1~q ),
	.datab(!\ic_fill_dp_offset_nxt[0]~1_combout ),
	.datac(!\ic_fill_dp_offset_nxt[1]~2_combout ),
	.datad(!\ic_fill_dp_offset_nxt[2]~0_combout ),
	.datae(!\ic_fill_valid_bits[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_fill_valid_bits_nxt~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_fill_valid_bits_nxt~4 .extended_lut = "off";
defparam \ic_fill_valid_bits_nxt~4 .lut_mask = 64'hFFFBFFFFFFFBFFFF;
defparam \ic_fill_valid_bits_nxt~4 .shared_arith = "off";

cyclonev_lcell_comb \ic_fill_valid_bits_nxt~5 (
	.dataa(!\D_ic_fill_starting_d1~q ),
	.datab(!\ic_fill_dp_offset_nxt[0]~1_combout ),
	.datac(!\ic_fill_dp_offset_nxt[1]~2_combout ),
	.datad(!\ic_fill_dp_offset_nxt[2]~0_combout ),
	.datae(!\ic_fill_valid_bits[3]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_fill_valid_bits_nxt~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_fill_valid_bits_nxt~5 .extended_lut = "off";
defparam \ic_fill_valid_bits_nxt~5 .lut_mask = 64'hFFBFFFFFFFBFFFFF;
defparam \ic_fill_valid_bits_nxt~5 .shared_arith = "off";

cyclonev_lcell_comb \ic_fill_valid_bits_nxt~6 (
	.dataa(!\D_ic_fill_starting_d1~q ),
	.datab(!\ic_fill_dp_offset_nxt[0]~1_combout ),
	.datac(!\ic_fill_dp_offset_nxt[1]~2_combout ),
	.datad(!\ic_fill_dp_offset_nxt[2]~0_combout ),
	.datae(!\ic_fill_valid_bits[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_fill_valid_bits_nxt~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_fill_valid_bits_nxt~6 .extended_lut = "off";
defparam \ic_fill_valid_bits_nxt~6 .lut_mask = 64'hFFFEFFFFFFFEFFFF;
defparam \ic_fill_valid_bits_nxt~6 .shared_arith = "off";

cyclonev_lcell_comb \ic_fill_valid_bits_nxt~7 (
	.dataa(!\D_ic_fill_starting_d1~q ),
	.datab(!\ic_fill_dp_offset_nxt[0]~1_combout ),
	.datac(!\ic_fill_dp_offset_nxt[1]~2_combout ),
	.datad(!\ic_fill_dp_offset_nxt[2]~0_combout ),
	.datae(!\ic_fill_valid_bits[2]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_fill_valid_bits_nxt~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_fill_valid_bits_nxt~7 .extended_lut = "off";
defparam \ic_fill_valid_bits_nxt~7 .lut_mask = 64'hFFEFFFFFFFEFFFFF;
defparam \ic_fill_valid_bits_nxt~7 .shared_arith = "off";

cyclonev_lcell_comb \ic_tag_clr_valid_bits~0 (
	.dataa(!\ic_tag_clr_valid_bits_nxt~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_tag_clr_valid_bits~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_tag_clr_valid_bits~0 .extended_lut = "off";
defparam \ic_tag_clr_valid_bits~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \ic_tag_clr_valid_bits~0 .shared_arith = "off";

dffeas \M_st_data[8] (
	.clk(clk_clk),
	.d(\E_stb_data[0]~2_combout ),
	.asdata(\E_stw_data[8]~11_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Equal0~0_combout ),
	.ena(\W_stall~combout ),
	.q(M_st_data_8),
	.prn(vcc));
defparam \M_st_data[8] .is_wysiwyg = "true";
defparam \M_st_data[8] .power_up = "low";

dffeas \M_st_data[9] (
	.clk(clk_clk),
	.d(\E_stb_data[1]~12_combout ),
	.asdata(\E_stw_data[9]~12_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Equal0~0_combout ),
	.ena(\W_stall~combout ),
	.q(M_st_data_9),
	.prn(vcc));
defparam \M_st_data[9] .is_wysiwyg = "true";
defparam \M_st_data[9] .power_up = "low";

dffeas \M_st_data[16] (
	.clk(clk_clk),
	.d(\E_stb_data[0]~2_combout ),
	.asdata(\E_stw_data[16]~2_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_iw[4]~q ),
	.ena(\W_stall~combout ),
	.q(M_st_data_16),
	.prn(vcc));
defparam \M_st_data[16] .is_wysiwyg = "true";
defparam \M_st_data[16] .power_up = "low";

dffeas \M_st_data[21] (
	.clk(clk_clk),
	.d(\E_stb_data[5]~14_combout ),
	.asdata(\E_stw_data[21]~21_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_iw[4]~q ),
	.ena(\W_stall~combout ),
	.q(M_st_data_21),
	.prn(vcc));
defparam \M_st_data[21] .is_wysiwyg = "true";
defparam \M_st_data[21] .power_up = "low";

dffeas \M_st_data[13] (
	.clk(clk_clk),
	.d(\E_stb_data[5]~14_combout ),
	.asdata(\E_stw_data[13]~13_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Equal0~0_combout ),
	.ena(\W_stall~combout ),
	.q(M_st_data_13),
	.prn(vcc));
defparam \M_st_data[13] .is_wysiwyg = "true";
defparam \M_st_data[13] .power_up = "low";

dffeas \M_st_data[20] (
	.clk(clk_clk),
	.d(\E_stb_data[4]~5_combout ),
	.asdata(\E_stw_data[20]~25_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_iw[4]~q ),
	.ena(\W_stall~combout ),
	.q(M_st_data_20),
	.prn(vcc));
defparam \M_st_data[20] .is_wysiwyg = "true";
defparam \M_st_data[20] .power_up = "low";

dffeas \M_st_data[12] (
	.clk(clk_clk),
	.d(\E_stb_data[4]~5_combout ),
	.asdata(\E_stw_data[12]~5_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Equal0~0_combout ),
	.ena(\W_stall~combout ),
	.q(M_st_data_12),
	.prn(vcc));
defparam \M_st_data[12] .is_wysiwyg = "true";
defparam \M_st_data[12] .power_up = "low";

dffeas \M_st_data[22] (
	.clk(clk_clk),
	.d(\E_stb_data[6]~8_combout ),
	.asdata(\E_stw_data[22]~31_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_iw[4]~q ),
	.ena(\W_stall~combout ),
	.q(M_st_data_22),
	.prn(vcc));
defparam \M_st_data[22] .is_wysiwyg = "true";
defparam \M_st_data[22] .power_up = "low";

dffeas \M_st_data[14] (
	.clk(clk_clk),
	.d(\E_stb_data[6]~8_combout ),
	.asdata(\E_stw_data[14]~4_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Equal0~0_combout ),
	.ena(\W_stall~combout ),
	.q(M_st_data_14),
	.prn(vcc));
defparam \M_st_data[14] .is_wysiwyg = "true";
defparam \M_st_data[14] .power_up = "low";

dffeas \M_st_data[23] (
	.clk(clk_clk),
	.d(\E_stb_data[7]~15_combout ),
	.asdata(\E_stw_data[23]~36_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_iw[4]~q ),
	.ena(\W_stall~combout ),
	.q(M_st_data_23),
	.prn(vcc));
defparam \M_st_data[23] .is_wysiwyg = "true";
defparam \M_st_data[23] .power_up = "low";

dffeas \M_st_data[15] (
	.clk(clk_clk),
	.d(\E_stb_data[7]~15_combout ),
	.asdata(\E_stw_data[15]~3_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Equal0~0_combout ),
	.ena(\W_stall~combout ),
	.q(M_st_data_15),
	.prn(vcc));
defparam \M_st_data[15] .is_wysiwyg = "true";
defparam \M_st_data[15] .power_up = "low";

dffeas \M_st_data[11] (
	.clk(clk_clk),
	.d(\E_stb_data[3]~13_combout ),
	.asdata(\E_stw_data[11]~14_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Equal0~0_combout ),
	.ena(\W_stall~combout ),
	.q(M_st_data_11),
	.prn(vcc));
defparam \M_st_data[11] .is_wysiwyg = "true";
defparam \M_st_data[11] .power_up = "low";

dffeas \M_st_data[10] (
	.clk(clk_clk),
	.d(\E_stb_data[2]~11_combout ),
	.asdata(\E_stw_data[10]~8_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Equal0~0_combout ),
	.ena(\W_stall~combout ),
	.q(M_st_data_10),
	.prn(vcc));
defparam \M_st_data[10] .is_wysiwyg = "true";
defparam \M_st_data[10] .power_up = "low";

dffeas \M_st_data[19] (
	.clk(clk_clk),
	.d(\E_stb_data[3]~13_combout ),
	.asdata(\E_stw_data[19]~42_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_iw[4]~q ),
	.ena(\W_stall~combout ),
	.q(M_st_data_19),
	.prn(vcc));
defparam \M_st_data[19] .is_wysiwyg = "true";
defparam \M_st_data[19] .power_up = "low";

dffeas \M_st_data[18] (
	.clk(clk_clk),
	.d(\E_stb_data[2]~11_combout ),
	.asdata(\E_stw_data[18]~34_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_iw[4]~q ),
	.ena(\W_stall~combout ),
	.q(M_st_data_18),
	.prn(vcc));
defparam \M_st_data[18] .is_wysiwyg = "true";
defparam \M_st_data[18] .power_up = "low";

dffeas \M_st_data[17] (
	.clk(clk_clk),
	.d(\E_stb_data[1]~12_combout ),
	.asdata(\E_stw_data[17]~35_combout ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_iw[4]~q ),
	.ena(\W_stall~combout ),
	.q(M_st_data_17),
	.prn(vcc));
defparam \M_st_data[17] .is_wysiwyg = "true";
defparam \M_st_data[17] .power_up = "low";

dffeas \M_st_data[0] (
	.clk(clk_clk),
	.d(\E_stb_data[0]~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(M_st_data_0),
	.prn(vcc));
defparam \M_st_data[0] .is_wysiwyg = "true";
defparam \M_st_data[0] .power_up = "low";

dffeas clr_break_line(
	.clk(clk_clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(clr_break_line1),
	.prn(vcc));
defparam clr_break_line.is_wysiwyg = "true";
defparam clr_break_line.power_up = "low";

dffeas d_write(
	.clk(clk_clk),
	.d(\d_write_nxt~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_write1),
	.prn(vcc));
defparam d_write.is_wysiwyg = "true";
defparam d_write.power_up = "low";

dffeas \M_alu_result[5] (
	.clk(clk_clk),
	.d(\E_alu_result[5]~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(M_alu_result_5),
	.prn(vcc));
defparam \M_alu_result[5] .is_wysiwyg = "true";
defparam \M_alu_result[5] .power_up = "low";

dffeas \M_alu_result[4] (
	.clk(clk_clk),
	.d(\E_alu_result[4]~4_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(M_alu_result_4),
	.prn(vcc));
defparam \M_alu_result[4] .is_wysiwyg = "true";
defparam \M_alu_result[4] .power_up = "low";

dffeas \M_alu_result[6] (
	.clk(clk_clk),
	.d(\E_alu_result[6]~5_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(M_alu_result_6),
	.prn(vcc));
defparam \M_alu_result[6] .is_wysiwyg = "true";
defparam \M_alu_result[6] .power_up = "low";

dffeas \M_alu_result[16] (
	.clk(clk_clk),
	.d(\E_wrctl_data_ienable_reg_irq16~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(M_alu_result_16),
	.prn(vcc));
defparam \M_alu_result[16] .is_wysiwyg = "true";
defparam \M_alu_result[16] .power_up = "low";

dffeas \M_alu_result[15] (
	.clk(clk_clk),
	.d(\E_alu_result[15]~7_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(M_alu_result_15),
	.prn(vcc));
defparam \M_alu_result[15] .is_wysiwyg = "true";
defparam \M_alu_result[15] .power_up = "low";

dffeas \M_alu_result[14] (
	.clk(clk_clk),
	.d(\E_alu_result[14]~9_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(M_alu_result_14),
	.prn(vcc));
defparam \M_alu_result[14] .is_wysiwyg = "true";
defparam \M_alu_result[14] .power_up = "low";

dffeas \M_alu_result[13] (
	.clk(clk_clk),
	.d(\E_alu_result[13]~11_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(M_alu_result_13),
	.prn(vcc));
defparam \M_alu_result[13] .is_wysiwyg = "true";
defparam \M_alu_result[13] .power_up = "low";

dffeas \M_alu_result[12] (
	.clk(clk_clk),
	.d(\E_alu_result[12]~13_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(M_alu_result_12),
	.prn(vcc));
defparam \M_alu_result[12] .is_wysiwyg = "true";
defparam \M_alu_result[12] .power_up = "low";

dffeas \M_alu_result[11] (
	.clk(clk_clk),
	.d(\E_alu_result[11]~15_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(M_alu_result_11),
	.prn(vcc));
defparam \M_alu_result[11] .is_wysiwyg = "true";
defparam \M_alu_result[11] .power_up = "low";

dffeas \M_alu_result[10] (
	.clk(clk_clk),
	.d(\E_alu_result[10]~16_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(M_alu_result_10),
	.prn(vcc));
defparam \M_alu_result[10] .is_wysiwyg = "true";
defparam \M_alu_result[10] .power_up = "low";

dffeas \M_alu_result[9] (
	.clk(clk_clk),
	.d(\E_alu_result[9]~18_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(M_alu_result_9),
	.prn(vcc));
defparam \M_alu_result[9] .is_wysiwyg = "true";
defparam \M_alu_result[9] .power_up = "low";

dffeas \M_alu_result[8] (
	.clk(clk_clk),
	.d(\E_alu_result[8]~19_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(M_alu_result_8),
	.prn(vcc));
defparam \M_alu_result[8] .is_wysiwyg = "true";
defparam \M_alu_result[8] .power_up = "low";

dffeas \M_alu_result[7] (
	.clk(clk_clk),
	.d(\E_alu_result[7]~21_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(M_alu_result_7),
	.prn(vcc));
defparam \M_alu_result[7] .is_wysiwyg = "true";
defparam \M_alu_result[7] .power_up = "low";

dffeas \M_alu_result[3] (
	.clk(clk_clk),
	.d(\E_alu_result[3]~23_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(M_alu_result_3),
	.prn(vcc));
defparam \M_alu_result[3] .is_wysiwyg = "true";
defparam \M_alu_result[3] .power_up = "low";

dffeas \M_alu_result[2] (
	.clk(clk_clk),
	.d(\E_alu_result[2]~25_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(M_alu_result_2),
	.prn(vcc));
defparam \M_alu_result[2] .is_wysiwyg = "true";
defparam \M_alu_result[2] .power_up = "low";

dffeas \M_st_data[1] (
	.clk(clk_clk),
	.d(\E_stb_data[1]~12_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(M_st_data_1),
	.prn(vcc));
defparam \M_st_data[1] .is_wysiwyg = "true";
defparam \M_st_data[1] .power_up = "low";

dffeas \M_st_data[2] (
	.clk(clk_clk),
	.d(\E_stb_data[2]~11_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(M_st_data_2),
	.prn(vcc));
defparam \M_st_data[2] .is_wysiwyg = "true";
defparam \M_st_data[2] .power_up = "low";

dffeas \M_st_data[3] (
	.clk(clk_clk),
	.d(\E_stb_data[3]~13_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(M_st_data_3),
	.prn(vcc));
defparam \M_st_data[3] .is_wysiwyg = "true";
defparam \M_st_data[3] .power_up = "low";

dffeas \M_st_data[4] (
	.clk(clk_clk),
	.d(\E_stb_data[4]~5_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(M_st_data_4),
	.prn(vcc));
defparam \M_st_data[4] .is_wysiwyg = "true";
defparam \M_st_data[4] .power_up = "low";

dffeas \M_st_data[5] (
	.clk(clk_clk),
	.d(\E_stb_data[5]~14_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(M_st_data_5),
	.prn(vcc));
defparam \M_st_data[5] .is_wysiwyg = "true";
defparam \M_st_data[5] .power_up = "low";

dffeas \M_st_data[6] (
	.clk(clk_clk),
	.d(\E_stb_data[6]~8_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(M_st_data_6),
	.prn(vcc));
defparam \M_st_data[6] .is_wysiwyg = "true";
defparam \M_st_data[6] .power_up = "low";

dffeas \M_st_data[7] (
	.clk(clk_clk),
	.d(\E_stb_data[7]~15_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(M_st_data_7),
	.prn(vcc));
defparam \M_st_data[7] .is_wysiwyg = "true";
defparam \M_st_data[7] .power_up = "low";

dffeas d_read(
	.clk(clk_clk),
	.d(\d_read_nxt~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_read1),
	.prn(vcc));
defparam d_read.is_wysiwyg = "true";
defparam d_read.power_up = "low";

dffeas hbreak_enabled(
	.clk(clk_clk),
	.d(\hbreak_enabled~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(hbreak_enabled1),
	.prn(vcc));
defparam hbreak_enabled.is_wysiwyg = "true";
defparam hbreak_enabled.power_up = "low";

dffeas i_read(
	.clk(clk_clk),
	.d(\i_read_nxt~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(i_read1),
	.prn(vcc));
defparam i_read.is_wysiwyg = "true";
defparam i_read.power_up = "low";

dffeas \ic_fill_tag[5] (
	.clk(clk_clk),
	.d(\D_pc[14]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\D_ic_fill_starting~0_combout ),
	.q(ic_fill_tag_5),
	.prn(vcc));
defparam \ic_fill_tag[5] .is_wysiwyg = "true";
defparam \ic_fill_tag[5] .power_up = "low";

dffeas \ic_fill_tag[4] (
	.clk(clk_clk),
	.d(\D_pc[13]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\D_ic_fill_starting~0_combout ),
	.q(ic_fill_tag_4),
	.prn(vcc));
defparam \ic_fill_tag[4] .is_wysiwyg = "true";
defparam \ic_fill_tag[4] .power_up = "low";

dffeas \ic_fill_tag[3] (
	.clk(clk_clk),
	.d(\D_pc[12]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\D_ic_fill_starting~0_combout ),
	.q(ic_fill_tag_3),
	.prn(vcc));
defparam \ic_fill_tag[3] .is_wysiwyg = "true";
defparam \ic_fill_tag[3] .power_up = "low";

dffeas \ic_fill_tag[2] (
	.clk(clk_clk),
	.d(\D_pc[11]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\D_ic_fill_starting~0_combout ),
	.q(ic_fill_tag_2),
	.prn(vcc));
defparam \ic_fill_tag[2] .is_wysiwyg = "true";
defparam \ic_fill_tag[2] .power_up = "low";

dffeas \ic_fill_tag[1] (
	.clk(clk_clk),
	.d(\D_pc[10]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\D_ic_fill_starting~0_combout ),
	.q(ic_fill_tag_1),
	.prn(vcc));
defparam \ic_fill_tag[1] .is_wysiwyg = "true";
defparam \ic_fill_tag[1] .power_up = "low";

dffeas \ic_fill_tag[0] (
	.clk(clk_clk),
	.d(\D_pc[9]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\D_ic_fill_starting~0_combout ),
	.q(ic_fill_tag_0),
	.prn(vcc));
defparam \ic_fill_tag[0] .is_wysiwyg = "true";
defparam \ic_fill_tag[0] .power_up = "low";

dffeas \ic_fill_line[5] (
	.clk(clk_clk),
	.d(\ic_tag_wraddress_nxt~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(ic_fill_line_5),
	.prn(vcc));
defparam \ic_fill_line[5] .is_wysiwyg = "true";
defparam \ic_fill_line[5] .power_up = "low";

dffeas \ic_fill_line[0] (
	.clk(clk_clk),
	.d(\ic_tag_wraddress_nxt~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(ic_fill_line_0),
	.prn(vcc));
defparam \ic_fill_line[0] .is_wysiwyg = "true";
defparam \ic_fill_line[0] .power_up = "low";

dffeas \ic_fill_line[1] (
	.clk(clk_clk),
	.d(\ic_tag_wraddress_nxt~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(ic_fill_line_1),
	.prn(vcc));
defparam \ic_fill_line[1] .is_wysiwyg = "true";
defparam \ic_fill_line[1] .power_up = "low";

dffeas \ic_fill_line[2] (
	.clk(clk_clk),
	.d(\ic_tag_wraddress_nxt~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(ic_fill_line_2),
	.prn(vcc));
defparam \ic_fill_line[2] .is_wysiwyg = "true";
defparam \ic_fill_line[2] .power_up = "low";

dffeas \ic_fill_line[3] (
	.clk(clk_clk),
	.d(\ic_tag_wraddress_nxt~4_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(ic_fill_line_3),
	.prn(vcc));
defparam \ic_fill_line[3] .is_wysiwyg = "true";
defparam \ic_fill_line[3] .power_up = "low";

dffeas \ic_fill_line[4] (
	.clk(clk_clk),
	.d(\ic_tag_wraddress_nxt~5_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(ic_fill_line_4),
	.prn(vcc));
defparam \ic_fill_line[4] .is_wysiwyg = "true";
defparam \ic_fill_line[4] .power_up = "low";

dffeas \ic_fill_ap_offset[0] (
	.clk(clk_clk),
	.d(\ic_fill_ap_offset_nxt[0]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ic_fill_ap_cnt[2]~0_combout ),
	.q(ic_fill_ap_offset_0),
	.prn(vcc));
defparam \ic_fill_ap_offset[0] .is_wysiwyg = "true";
defparam \ic_fill_ap_offset[0] .power_up = "low";

dffeas \ic_fill_ap_offset[1] (
	.clk(clk_clk),
	.d(\ic_fill_ap_offset_nxt[1]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ic_fill_ap_cnt[2]~0_combout ),
	.q(ic_fill_ap_offset_1),
	.prn(vcc));
defparam \ic_fill_ap_offset[1] .is_wysiwyg = "true";
defparam \ic_fill_ap_offset[1] .power_up = "low";

dffeas \ic_fill_ap_offset[2] (
	.clk(clk_clk),
	.d(\ic_fill_ap_offset_nxt[2]~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ic_fill_ap_cnt[2]~0_combout ),
	.q(ic_fill_ap_offset_2),
	.prn(vcc));
defparam \ic_fill_ap_offset[2] .is_wysiwyg = "true";
defparam \ic_fill_ap_offset[2] .power_up = "low";

dffeas \M_mem_byte_en[0] (
	.clk(clk_clk),
	.d(\E_mem_byte_en~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(M_mem_byte_en_0),
	.prn(vcc));
defparam \M_mem_byte_en[0] .is_wysiwyg = "true";
defparam \M_mem_byte_en[0] .power_up = "low";

dffeas \M_mem_byte_en[2] (
	.clk(clk_clk),
	.d(\E_mem_byte_en[2]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(M_mem_byte_en_2),
	.prn(vcc));
defparam \M_mem_byte_en[2] .is_wysiwyg = "true";
defparam \M_mem_byte_en[2] .power_up = "low";

dffeas \M_mem_byte_en[1] (
	.clk(clk_clk),
	.d(\E_mem_byte_en[1]~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(M_mem_byte_en_1),
	.prn(vcc));
defparam \M_mem_byte_en[1] .is_wysiwyg = "true";
defparam \M_mem_byte_en[1] .power_up = "low";

dffeas \M_st_data[24] (
	.clk(clk_clk),
	.d(\E_st_data[24]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(M_st_data_24),
	.prn(vcc));
defparam \M_st_data[24] .is_wysiwyg = "true";
defparam \M_st_data[24] .power_up = "low";

dffeas \M_mem_byte_en[3] (
	.clk(clk_clk),
	.d(\E_mem_byte_en[3]~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(M_mem_byte_en_3),
	.prn(vcc));
defparam \M_mem_byte_en[3] .is_wysiwyg = "true";
defparam \M_mem_byte_en[3] .power_up = "low";

dffeas \M_st_data[29] (
	.clk(clk_clk),
	.d(\E_st_data[29]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(M_st_data_29),
	.prn(vcc));
defparam \M_st_data[29] .is_wysiwyg = "true";
defparam \M_st_data[29] .power_up = "low";

dffeas \M_st_data[28] (
	.clk(clk_clk),
	.d(\E_st_data[28]~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(M_st_data_28),
	.prn(vcc));
defparam \M_st_data[28] .is_wysiwyg = "true";
defparam \M_st_data[28] .power_up = "low";

dffeas \M_st_data[30] (
	.clk(clk_clk),
	.d(\E_st_data[30]~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(M_st_data_30),
	.prn(vcc));
defparam \M_st_data[30] .is_wysiwyg = "true";
defparam \M_st_data[30] .power_up = "low";

dffeas \M_st_data[31] (
	.clk(clk_clk),
	.d(\E_st_data[31]~5_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(M_st_data_31),
	.prn(vcc));
defparam \M_st_data[31] .is_wysiwyg = "true";
defparam \M_st_data[31] .power_up = "low";

dffeas \M_st_data[27] (
	.clk(clk_clk),
	.d(\E_st_data[27]~6_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(M_st_data_27),
	.prn(vcc));
defparam \M_st_data[27] .is_wysiwyg = "true";
defparam \M_st_data[27] .power_up = "low";

dffeas \M_st_data[26] (
	.clk(clk_clk),
	.d(\E_st_data[26]~7_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(M_st_data_26),
	.prn(vcc));
defparam \M_st_data[26] .is_wysiwyg = "true";
defparam \M_st_data[26] .power_up = "low";

dffeas \M_st_data[25] (
	.clk(clk_clk),
	.d(\E_st_data[25]~8_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(M_st_data_25),
	.prn(vcc));
defparam \M_st_data[25] .is_wysiwyg = "true";
defparam \M_st_data[25] .power_up = "low";

cyclonev_lcell_comb \F_iw[0]~2 (
	.dataa(!\intr_req~0_combout ),
	.datab(!\processor_cpu_ic_data|the_altsyncram|auto_generated|q_b[0] ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[0]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[0]~2 .extended_lut = "off";
defparam \F_iw[0]~2 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \F_iw[0]~2 .shared_arith = "off";

cyclonev_lcell_comb \F_iw[14]~12 (
	.dataa(!\intr_req~0_combout ),
	.datab(!\processor_cpu_ic_data|the_altsyncram|auto_generated|q_b[14] ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[14]~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[14]~12 .extended_lut = "off";
defparam \F_iw[14]~12 .lut_mask = 64'h7777777777777777;
defparam \F_iw[14]~12 .shared_arith = "off";

cyclonev_lcell_comb \av_ld_data_transfer~0 (
	.dataa(!d_read1),
	.datab(!WideOr1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_ld_data_transfer~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_ld_data_transfer~0 .extended_lut = "off";
defparam \av_ld_data_transfer~0 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \av_ld_data_transfer~0 .shared_arith = "off";

dffeas av_ld_aligning_data(
	.clk(clk_clk),
	.d(\av_ld_data_transfer~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\av_ld_aligning_data~q ),
	.prn(vcc));
defparam av_ld_aligning_data.is_wysiwyg = "true";
defparam av_ld_aligning_data.power_up = "low";

dffeas av_ld_or_div_done(
	.clk(clk_clk),
	.d(\av_ld_aligning_data~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\av_ld_or_div_done~q ),
	.prn(vcc));
defparam av_ld_or_div_done.is_wysiwyg = "true";
defparam av_ld_or_div_done.power_up = "low";

cyclonev_lcell_comb \F_iw[5]~7 (
	.dataa(!\F_iw~1_combout ),
	.datab(!\intr_req~0_combout ),
	.datac(!\processor_cpu_ic_data|the_altsyncram|auto_generated|q_b[5] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[5]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[5]~7 .extended_lut = "off";
defparam \F_iw[5]~7 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \F_iw[5]~7 .shared_arith = "off";

dffeas \D_iw[5] (
	.clk(clk_clk),
	.d(\F_iw[5]~7_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\D_iw[5]~q ),
	.prn(vcc));
defparam \D_iw[5] .is_wysiwyg = "true";
defparam \D_iw[5] .power_up = "low";

dffeas \E_iw[5] (
	.clk(clk_clk),
	.d(\D_iw[5]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_iw[5]~q ),
	.prn(vcc));
defparam \E_iw[5] .is_wysiwyg = "true";
defparam \E_iw[5] .power_up = "low";

cyclonev_lcell_comb \F_iw[4]~6 (
	.dataa(!\F_iw~1_combout ),
	.datab(!\intr_req~0_combout ),
	.datac(!\processor_cpu_ic_data|the_altsyncram|auto_generated|q_b[4] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[4]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[4]~6 .extended_lut = "off";
defparam \F_iw[4]~6 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \F_iw[4]~6 .shared_arith = "off";

dffeas \D_iw[4] (
	.clk(clk_clk),
	.d(\F_iw[4]~6_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\D_iw[4]~q ),
	.prn(vcc));
defparam \D_iw[4] .is_wysiwyg = "true";
defparam \D_iw[4] .power_up = "low";

dffeas \E_iw[4] (
	.clk(clk_clk),
	.d(\D_iw[4]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_iw[4]~q ),
	.prn(vcc));
defparam \E_iw[4] .is_wysiwyg = "true";
defparam \E_iw[4] .power_up = "low";

cyclonev_lcell_comb \F_iw[3]~5 (
	.dataa(!\F_iw~1_combout ),
	.datab(!\intr_req~0_combout ),
	.datac(!\processor_cpu_ic_data|the_altsyncram|auto_generated|q_b[3] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[3]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[3]~5 .extended_lut = "off";
defparam \F_iw[3]~5 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \F_iw[3]~5 .shared_arith = "off";

dffeas \D_iw[3] (
	.clk(clk_clk),
	.d(\F_iw[3]~5_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\D_iw[3]~q ),
	.prn(vcc));
defparam \D_iw[3] .is_wysiwyg = "true";
defparam \D_iw[3] .power_up = "low";

dffeas \E_iw[3] (
	.clk(clk_clk),
	.d(\D_iw[3]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_iw[3]~q ),
	.prn(vcc));
defparam \E_iw[3] .is_wysiwyg = "true";
defparam \E_iw[3] .power_up = "low";

cyclonev_lcell_comb \F_iw[2]~4 (
	.dataa(!\intr_req~0_combout ),
	.datab(!\processor_cpu_ic_data|the_altsyncram|auto_generated|q_b[2] ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[2]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[2]~4 .extended_lut = "off";
defparam \F_iw[2]~4 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \F_iw[2]~4 .shared_arith = "off";

dffeas \D_iw[2] (
	.clk(clk_clk),
	.d(\F_iw[2]~4_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\F_iw~1_combout ),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\D_iw[2]~q ),
	.prn(vcc));
defparam \D_iw[2] .is_wysiwyg = "true";
defparam \D_iw[2] .power_up = "low";

dffeas \E_iw[2] (
	.clk(clk_clk),
	.d(\D_iw[2]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_iw[2]~q ),
	.prn(vcc));
defparam \E_iw[2] .is_wysiwyg = "true";
defparam \E_iw[2] .power_up = "low";

cyclonev_lcell_comb \F_iw[1]~3 (
	.dataa(!\F_iw~1_combout ),
	.datab(!\intr_req~0_combout ),
	.datac(!\processor_cpu_ic_data|the_altsyncram|auto_generated|q_b[1] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[1]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[1]~3 .extended_lut = "off";
defparam \F_iw[1]~3 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \F_iw[1]~3 .shared_arith = "off";

dffeas \D_iw[1] (
	.clk(clk_clk),
	.d(\F_iw[1]~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\D_iw[1]~q ),
	.prn(vcc));
defparam \D_iw[1] .is_wysiwyg = "true";
defparam \D_iw[1] .power_up = "low";

dffeas \E_iw[1] (
	.clk(clk_clk),
	.d(\D_iw[1]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_iw[1]~q ),
	.prn(vcc));
defparam \E_iw[1] .is_wysiwyg = "true";
defparam \E_iw[1] .power_up = "low";

dffeas \E_iw[0] (
	.clk(clk_clk),
	.d(\D_iw[0]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_iw[0]~q ),
	.prn(vcc));
defparam \E_iw[0] .is_wysiwyg = "true";
defparam \E_iw[0] .power_up = "low";

cyclonev_lcell_comb \Equal130~0 (
	.dataa(!\E_iw[5]~q ),
	.datab(!\E_iw[4]~q ),
	.datac(!\E_iw[3]~q ),
	.datad(!\E_iw[2]~q ),
	.datae(!\E_iw[1]~q ),
	.dataf(!\E_iw[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal130~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal130~0 .extended_lut = "off";
defparam \Equal130~0 .lut_mask = 64'hFFFFFFFFFF7FFFFF;
defparam \Equal130~0 .shared_arith = "off";

cyclonev_lcell_comb \F_iw[12]~13 (
	.dataa(!\intr_req~0_combout ),
	.datab(!\processor_cpu_ic_data|the_altsyncram|auto_generated|q_b[12] ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[12]~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[12]~13 .extended_lut = "off";
defparam \F_iw[12]~13 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \F_iw[12]~13 .shared_arith = "off";

dffeas \D_iw[12] (
	.clk(clk_clk),
	.d(\F_iw[12]~13_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\F_iw~1_combout ),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\D_iw[12]~q ),
	.prn(vcc));
defparam \D_iw[12] .is_wysiwyg = "true";
defparam \D_iw[12] .power_up = "low";

dffeas \E_iw[12] (
	.clk(clk_clk),
	.d(\D_iw[12]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_iw[12]~q ),
	.prn(vcc));
defparam \E_iw[12] .is_wysiwyg = "true";
defparam \E_iw[12] .power_up = "low";

cyclonev_lcell_comb \F_iw[11]~14 (
	.dataa(!\F_iw~1_combout ),
	.datab(!\intr_req~0_combout ),
	.datac(!\processor_cpu_ic_data|the_altsyncram|auto_generated|q_b[11] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[11]~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[11]~14 .extended_lut = "off";
defparam \F_iw[11]~14 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \F_iw[11]~14 .shared_arith = "off";

dffeas \D_iw[11] (
	.clk(clk_clk),
	.d(\F_iw[11]~14_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\D_iw[11]~q ),
	.prn(vcc));
defparam \D_iw[11] .is_wysiwyg = "true";
defparam \D_iw[11] .power_up = "low";

dffeas \E_iw[11] (
	.clk(clk_clk),
	.d(\D_iw[11]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_iw[11]~q ),
	.prn(vcc));
defparam \E_iw[11] .is_wysiwyg = "true";
defparam \E_iw[11] .power_up = "low";

cyclonev_lcell_comb \E_op_eret~0 (
	.dataa(!\E_iw[12]~q ),
	.datab(!\E_iw[11]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_op_eret~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_op_eret~0 .extended_lut = "off";
defparam \E_op_eret~0 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \E_op_eret~0 .shared_arith = "off";

cyclonev_lcell_comb \F_iw[16]~15 (
	.dataa(!\F_iw~1_combout ),
	.datab(!\intr_req~0_combout ),
	.datac(!\processor_cpu_ic_data|the_altsyncram|auto_generated|q_b[16] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[16]~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[16]~15 .extended_lut = "off";
defparam \F_iw[16]~15 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \F_iw[16]~15 .shared_arith = "off";

dffeas \D_iw[16] (
	.clk(clk_clk),
	.d(\F_iw[16]~15_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\D_iw[16]~q ),
	.prn(vcc));
defparam \D_iw[16] .is_wysiwyg = "true";
defparam \D_iw[16] .power_up = "low";

dffeas \E_iw[16] (
	.clk(clk_clk),
	.d(\D_iw[16]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_iw[16]~q ),
	.prn(vcc));
defparam \E_iw[16] .is_wysiwyg = "true";
defparam \E_iw[16] .power_up = "low";

cyclonev_lcell_comb \F_iw[15]~16 (
	.dataa(!\F_iw~1_combout ),
	.datab(!\intr_req~0_combout ),
	.datac(!\processor_cpu_ic_data|the_altsyncram|auto_generated|q_b[15] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[15]~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[15]~16 .extended_lut = "off";
defparam \F_iw[15]~16 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \F_iw[15]~16 .shared_arith = "off";

dffeas \D_iw[15] (
	.clk(clk_clk),
	.d(\F_iw[15]~16_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\D_iw[15]~q ),
	.prn(vcc));
defparam \D_iw[15] .is_wysiwyg = "true";
defparam \D_iw[15] .power_up = "low";

dffeas \E_iw[15] (
	.clk(clk_clk),
	.d(\D_iw[15]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_iw[15]~q ),
	.prn(vcc));
defparam \E_iw[15] .is_wysiwyg = "true";
defparam \E_iw[15] .power_up = "low";

cyclonev_lcell_comb \F_iw[13]~17 (
	.dataa(!\F_iw~1_combout ),
	.datab(!\intr_req~0_combout ),
	.datac(!\processor_cpu_ic_data|the_altsyncram|auto_generated|q_b[13] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[13]~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[13]~17 .extended_lut = "off";
defparam \F_iw[13]~17 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \F_iw[13]~17 .shared_arith = "off";

dffeas \D_iw[13] (
	.clk(clk_clk),
	.d(\F_iw[13]~17_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\D_iw[13]~q ),
	.prn(vcc));
defparam \D_iw[13] .is_wysiwyg = "true";
defparam \D_iw[13] .power_up = "low";

dffeas \E_iw[13] (
	.clk(clk_clk),
	.d(\D_iw[13]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_iw[13]~q ),
	.prn(vcc));
defparam \E_iw[13] .is_wysiwyg = "true";
defparam \E_iw[13] .power_up = "low";

cyclonev_lcell_comb \E_hbreak_req~0 (
	.dataa(!\E_iw[16]~q ),
	.datab(!\E_iw[15]~q ),
	.datac(!\E_iw[13]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_hbreak_req~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_hbreak_req~0 .extended_lut = "off";
defparam \E_hbreak_req~0 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \E_hbreak_req~0 .shared_arith = "off";

cyclonev_lcell_comb \wait_for_one_post_bret_inst~0 (
	.dataa(!\E_valid~0_combout ),
	.datab(!hbreak_enabled1),
	.datac(!\wait_for_one_post_bret_inst~q ),
	.datad(!\W_stall~combout ),
	.datae(!\the_processor_cpu_nios2_oci|the_processor_cpu_nios2_avalon_reg|oci_single_step_mode~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_for_one_post_bret_inst~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_for_one_post_bret_inst~0 .extended_lut = "off";
defparam \wait_for_one_post_bret_inst~0 .lut_mask = 64'hFFBFFFFFFFBFFFFF;
defparam \wait_for_one_post_bret_inst~0 .shared_arith = "off";

dffeas wait_for_one_post_bret_inst(
	.clk(clk_clk),
	.d(\wait_for_one_post_bret_inst~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wait_for_one_post_bret_inst~q ),
	.prn(vcc));
defparam wait_for_one_post_bret_inst.is_wysiwyg = "true";
defparam wait_for_one_post_bret_inst.power_up = "low";

cyclonev_lcell_comb \hbreak_req~0 (
	.dataa(!hbreak_enabled1),
	.datab(!\wait_for_one_post_bret_inst~q ),
	.datac(!\latched_oci_tb_hbreak_req~q ),
	.datad(!\the_processor_cpu_nios2_oci|the_processor_cpu_nios2_oci_debug|jtag_break~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\hbreak_req~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \hbreak_req~0 .extended_lut = "off";
defparam \hbreak_req~0 .lut_mask = 64'hEFFFEFFFEFFFEFFF;
defparam \hbreak_req~0 .shared_arith = "off";

cyclonev_lcell_comb \E_valid~1 (
	.dataa(!\E_iw[14]~q ),
	.datab(!\E_valid~0_combout ),
	.datac(!\Equal130~0_combout ),
	.datad(!\E_op_eret~0_combout ),
	.datae(!\E_hbreak_req~0_combout ),
	.dataf(!\hbreak_req~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_valid~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_valid~1 .extended_lut = "off";
defparam \E_valid~1 .lut_mask = 64'hFFFFFFFFBFFFFFFF;
defparam \E_valid~1 .shared_arith = "off";

dffeas M_valid_from_E(
	.clk(clk_clk),
	.d(\E_valid~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\M_valid_from_E~q ),
	.prn(vcc));
defparam M_valid_from_E.is_wysiwyg = "true";
defparam M_valid_from_E.power_up = "low";

cyclonev_lcell_comb \D_ctrl_ld~0 (
	.dataa(!\D_iw[4]~q ),
	.datab(!\D_iw[2]~q ),
	.datac(!\D_iw[1]~q ),
	.datad(!\D_iw[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_ld~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_ld~0 .extended_lut = "off";
defparam \D_ctrl_ld~0 .lut_mask = 64'hBFFFBFFFBFFFBFFF;
defparam \D_ctrl_ld~0 .shared_arith = "off";

dffeas E_ctrl_ld(
	.clk(clk_clk),
	.d(\D_ctrl_ld~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_ctrl_ld~q ),
	.prn(vcc));
defparam E_ctrl_ld.is_wysiwyg = "true";
defparam E_ctrl_ld.power_up = "low";

dffeas M_ctrl_ld(
	.clk(clk_clk),
	.d(\E_ctrl_ld~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\M_ctrl_ld~q ),
	.prn(vcc));
defparam M_ctrl_ld.is_wysiwyg = "true";
defparam M_ctrl_ld.power_up = "low";

cyclonev_lcell_comb \M_status_reg_pie~0 (
	.dataa(!d_write1),
	.datab(!d_read1),
	.datac(!WideOr1),
	.datad(!read_accepted),
	.datae(!\E_valid~1_combout ),
	.dataf(!\W_stall~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_status_reg_pie~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_status_reg_pie~0 .extended_lut = "off";
defparam \M_status_reg_pie~0 .lut_mask = 64'hB8FFFFFFFFFFFFFF;
defparam \M_status_reg_pie~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal4~0 (
	.dataa(!\D_iw[0]~q ),
	.datab(!\D_iw[1]~q ),
	.datac(!\D_iw[2]~q ),
	.datad(!\D_iw[3]~q ),
	.datae(!\D_iw[4]~q ),
	.dataf(!\D_iw[5]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal4~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal4~0 .extended_lut = "off";
defparam \Equal4~0 .lut_mask = 64'hFBFFFFFFFFFFFFFF;
defparam \Equal4~0 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_shift_logical~0 (
	.dataa(!\D_iw[12]~q ),
	.datab(!\D_iw[13]~q ),
	.datac(!\Equal4~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_shift_logical~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_shift_logical~0 .extended_lut = "off";
defparam \D_ctrl_shift_logical~0 .lut_mask = 64'hDFDFDFDFDFDFDFDF;
defparam \D_ctrl_shift_logical~0 .shared_arith = "off";

dffeas E_ctrl_shift_rot(
	.clk(clk_clk),
	.d(\D_ctrl_shift_logical~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_ctrl_shift_rot~q ),
	.prn(vcc));
defparam E_ctrl_shift_rot.is_wysiwyg = "true";
defparam E_ctrl_shift_rot.power_up = "low";

cyclonev_lcell_comb \D_ctrl_b_not_src~0 (
	.dataa(!\D_iw[5]~q ),
	.datab(!\D_iw[4]~q ),
	.datac(!\D_iw[3]~q ),
	.datad(!\D_iw[2]~q ),
	.datae(!\D_iw[1]~q ),
	.dataf(!\D_iw[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_b_not_src~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_b_not_src~0 .extended_lut = "off";
defparam \D_ctrl_b_not_src~0 .lut_mask = 64'hFDFFFFFFFFFFFDFF;
defparam \D_ctrl_b_not_src~0 .shared_arith = "off";

cyclonev_lcell_comb \D_wr_dst_reg~1 (
	.dataa(!\D_iw[2]~q ),
	.datab(!\D_iw[1]~q ),
	.datac(!\D_iw[0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_wr_dst_reg~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_wr_dst_reg~1 .extended_lut = "off";
defparam \D_wr_dst_reg~1 .lut_mask = 64'hDFDFDFDFDFDFDFDF;
defparam \D_wr_dst_reg~1 .shared_arith = "off";

cyclonev_lcell_comb D_ctrl_src2_choose_imm(
	.dataa(!\D_ctrl_b_not_src~0_combout ),
	.datab(!\D_iw[11]~q ),
	.datac(!\D_ctrl_shift_logical~0_combout ),
	.datad(!\D_wr_dst_reg~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_src2_choose_imm~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam D_ctrl_src2_choose_imm.extended_lut = "off";
defparam D_ctrl_src2_choose_imm.lut_mask = 64'hEFFFEFFFEFFFEFFF;
defparam D_ctrl_src2_choose_imm.shared_arith = "off";

dffeas E_ctrl_src2_choose_imm(
	.clk(clk_clk),
	.d(\D_ctrl_src2_choose_imm~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_ctrl_src2_choose_imm~q ),
	.prn(vcc));
defparam E_ctrl_src2_choose_imm.is_wysiwyg = "true";
defparam E_ctrl_src2_choose_imm.power_up = "low";

cyclonev_lcell_comb \F_iw[6]~25 (
	.dataa(!\intr_req~0_combout ),
	.datab(!\processor_cpu_ic_data|the_altsyncram|auto_generated|q_b[6] ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[6]~25_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[6]~25 .extended_lut = "off";
defparam \F_iw[6]~25 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \F_iw[6]~25 .shared_arith = "off";

dffeas \D_iw[6] (
	.clk(clk_clk),
	.d(\F_iw[6]~25_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\F_iw~1_combout ),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\D_iw[6]~q ),
	.prn(vcc));
defparam \D_iw[6] .is_wysiwyg = "true";
defparam \D_iw[6] .power_up = "low";

cyclonev_lcell_comb \D_ctrl_hi_imm16~0 (
	.dataa(!\D_iw[0]~q ),
	.datab(!\D_iw[1]~q ),
	.datac(!\D_iw[4]~q ),
	.datad(!\D_iw[3]~q ),
	.datae(!\D_iw[2]~q ),
	.dataf(!\D_iw[5]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_hi_imm16~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_hi_imm16~0 .extended_lut = "off";
defparam \D_ctrl_hi_imm16~0 .lut_mask = 64'hEFFFFFFFFFFFFFFF;
defparam \D_ctrl_hi_imm16~0 .shared_arith = "off";

dffeas \E_src2_imm[0] (
	.clk(clk_clk),
	.d(\D_iw[6]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\D_ctrl_hi_imm16~0_combout ),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_src2_imm[0]~q ),
	.prn(vcc));
defparam \E_src2_imm[0] .is_wysiwyg = "true";
defparam \E_src2_imm[0] .power_up = "low";

dffeas M_ctrl_shift_rot(
	.clk(clk_clk),
	.d(\E_ctrl_shift_rot~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\M_ctrl_shift_rot~q ),
	.prn(vcc));
defparam M_ctrl_shift_rot.is_wysiwyg = "true";
defparam M_ctrl_shift_rot.power_up = "low";

dffeas \d_readdata_d1[3] (
	.clk(clk_clk),
	.d(d_readdata[3]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d_readdata_d1[3]~q ),
	.prn(vcc));
defparam \d_readdata_d1[3] .is_wysiwyg = "true";
defparam \d_readdata_d1[3] .power_up = "low";

dffeas \d_readdata_d1[19] (
	.clk(clk_clk),
	.d(d_readdata[19]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d_readdata_d1[19]~q ),
	.prn(vcc));
defparam \d_readdata_d1[19] .is_wysiwyg = "true";
defparam \d_readdata_d1[19] .power_up = "low";

dffeas \d_readdata_d1[11] (
	.clk(clk_clk),
	.d(d_readdata[11]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d_readdata_d1[11]~q ),
	.prn(vcc));
defparam \d_readdata_d1[11] .is_wysiwyg = "true";
defparam \d_readdata_d1[11] .power_up = "low";

dffeas \d_readdata_d1[27] (
	.clk(clk_clk),
	.d(d_readdata[27]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d_readdata_d1[27]~q ),
	.prn(vcc));
defparam \d_readdata_d1[27] .is_wysiwyg = "true";
defparam \d_readdata_d1[27] .power_up = "low";

cyclonev_lcell_comb \D_ctrl_crst~0 (
	.dataa(!\D_iw[12]~q ),
	.datab(!\D_iw[13]~q ),
	.datac(!\Equal4~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_crst~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_crst~0 .extended_lut = "off";
defparam \D_ctrl_crst~0 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \D_ctrl_crst~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal107~1 (
	.dataa(!\D_iw[16]~q ),
	.datab(!\D_iw[15]~q ),
	.datac(!\D_iw[14]~q ),
	.datad(!\D_iw[11]~q ),
	.datae(!\D_ctrl_crst~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal107~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal107~1 .extended_lut = "off";
defparam \Equal107~1 .lut_mask = 64'hFFFDFFFFFFFDFFFF;
defparam \Equal107~1 .shared_arith = "off";

dffeas E_ctrl_rdctl_inst(
	.clk(clk_clk),
	.d(\Equal107~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_ctrl_rdctl_inst~q ),
	.prn(vcc));
defparam E_ctrl_rdctl_inst.is_wysiwyg = "true";
defparam E_ctrl_rdctl_inst.power_up = "low";

cyclonev_lcell_comb \D_ctrl_implicit_dst_retaddr~0 (
	.dataa(!\D_iw[0]~q ),
	.datab(!\D_iw[2]~q ),
	.datac(!\D_iw[3]~q ),
	.datad(!\D_iw[4]~q ),
	.datae(!\D_iw[5]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_implicit_dst_retaddr~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_implicit_dst_retaddr~0 .extended_lut = "off";
defparam \D_ctrl_implicit_dst_retaddr~0 .lut_mask = 64'hFFFFFFFEFFFFFFFE;
defparam \D_ctrl_implicit_dst_retaddr~0 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_retaddr~0 (
	.dataa(!\D_iw[16]~q ),
	.datab(!\D_iw[12]~q ),
	.datac(!\D_iw[15]~q ),
	.datad(!\D_iw[14]~q ),
	.datae(!\D_iw[11]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_retaddr~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_retaddr~0 .extended_lut = "off";
defparam \D_ctrl_retaddr~0 .lut_mask = 64'hEDDEFFFFEDDEFFFF;
defparam \D_ctrl_retaddr~0 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_break~0 (
	.dataa(!\D_iw[12]~q ),
	.datab(!\D_iw[15]~q ),
	.datac(!\D_iw[13]~q ),
	.datad(!\Equal4~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_break~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_break~0 .extended_lut = "off";
defparam \D_ctrl_break~0 .lut_mask = 64'hBFFFBFFFBFFFBFFF;
defparam \D_ctrl_break~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal4~1 (
	.dataa(!\D_iw[0]~q ),
	.datab(!\D_iw[1]~q ),
	.datac(!\D_iw[2]~q ),
	.datad(!\D_iw[3]~q ),
	.datae(!\D_iw[4]~q ),
	.dataf(!\D_iw[5]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal4~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal4~1 .extended_lut = "off";
defparam \Equal4~1 .lut_mask = 64'hFFFFFFEFFFFFFFFF;
defparam \Equal4~1 .shared_arith = "off";

cyclonev_lcell_comb \Equal107~0 (
	.dataa(!\D_iw[16]~q ),
	.datab(!\D_iw[12]~q ),
	.datac(!\D_iw[11]~q ),
	.datad(!\D_iw[13]~q ),
	.datae(!\Equal4~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal107~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal107~0 .extended_lut = "off";
defparam \Equal107~0 .lut_mask = 64'hBFFFFFFFBFFFFFFF;
defparam \Equal107~0 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_implicit_dst_eretaddr~0 (
	.dataa(!\D_iw[15]~q ),
	.datab(!\D_iw[14]~q ),
	.datac(!\Equal4~1_combout ),
	.datad(!\Equal107~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_implicit_dst_eretaddr~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_implicit_dst_eretaddr~0 .extended_lut = "off";
defparam \D_ctrl_implicit_dst_eretaddr~0 .lut_mask = 64'hFFFBFFFBFFFBFFFB;
defparam \D_ctrl_implicit_dst_eretaddr~0 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_exception~0 (
	.dataa(!\D_iw[16]~q ),
	.datab(!\D_iw[14]~q ),
	.datac(gnd),
	.datad(!\D_ctrl_break~0_combout ),
	.datae(!\D_ctrl_implicit_dst_eretaddr~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_exception~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_exception~0 .extended_lut = "off";
defparam \D_ctrl_exception~0 .lut_mask = 64'hFFEEFFFFFFEEFFFF;
defparam \D_ctrl_exception~0 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_retaddr~1 (
	.dataa(!\D_ctrl_implicit_dst_retaddr~0_combout ),
	.datab(!\D_ctrl_retaddr~0_combout ),
	.datac(!\D_iw[13]~q ),
	.datad(!\Equal4~0_combout ),
	.datae(!\D_ctrl_exception~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_retaddr~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_retaddr~1 .extended_lut = "off";
defparam \D_ctrl_retaddr~1 .lut_mask = 64'hFFFF7FFFFFFF7FFF;
defparam \D_ctrl_retaddr~1 .shared_arith = "off";

dffeas E_ctrl_retaddr(
	.clk(clk_clk),
	.d(\D_ctrl_retaddr~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_ctrl_retaddr~q ),
	.prn(vcc));
defparam E_ctrl_retaddr.is_wysiwyg = "true";
defparam E_ctrl_retaddr.power_up = "low";

cyclonev_lcell_comb \Equal4~5 (
	.dataa(!\D_iw[0]~q ),
	.datab(!\D_iw[1]~q ),
	.datac(!\D_iw[2]~q ),
	.datad(!\D_iw[3]~q ),
	.datae(!\D_iw[4]~q ),
	.dataf(!\D_iw[5]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal4~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal4~5 .extended_lut = "off";
defparam \Equal4~5 .lut_mask = 64'hFFFFFFFFFEFFFFFF;
defparam \Equal4~5 .shared_arith = "off";

cyclonev_lcell_comb \Equal4~6 (
	.dataa(!\D_iw[0]~q ),
	.datab(!\D_iw[1]~q ),
	.datac(!\D_iw[2]~q ),
	.datad(!\D_iw[3]~q ),
	.datae(!\D_iw[4]~q ),
	.dataf(!\D_iw[5]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal4~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal4~6 .extended_lut = "off";
defparam \Equal4~6 .lut_mask = 64'hFFFFFFFEFFFFFFFF;
defparam \Equal4~6 .shared_arith = "off";

cyclonev_lcell_comb \Equal4~7 (
	.dataa(!\D_iw[0]~q ),
	.datab(!\D_iw[1]~q ),
	.datac(!\D_iw[2]~q ),
	.datad(!\D_iw[3]~q ),
	.datae(!\D_iw[4]~q ),
	.dataf(!\D_iw[5]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal4~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal4~7 .extended_lut = "off";
defparam \Equal4~7 .lut_mask = 64'hFFFFFEFFFFFFFFFF;
defparam \Equal4~7 .shared_arith = "off";

cyclonev_lcell_comb \Equal4~8 (
	.dataa(!\D_iw[0]~q ),
	.datab(!\D_iw[1]~q ),
	.datac(!\D_iw[2]~q ),
	.datad(!\D_iw[3]~q ),
	.datae(!\D_iw[4]~q ),
	.dataf(!\D_iw[5]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal4~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal4~8 .extended_lut = "off";
defparam \Equal4~8 .lut_mask = 64'hFFFEFFFFFFFFFFFF;
defparam \Equal4~8 .shared_arith = "off";

cyclonev_lcell_comb \Equal4~9 (
	.dataa(!\D_iw[0]~q ),
	.datab(!\D_iw[1]~q ),
	.datac(!\D_iw[2]~q ),
	.datad(!\D_iw[3]~q ),
	.datae(!\D_iw[4]~q ),
	.dataf(!\D_iw[5]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal4~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal4~9 .extended_lut = "off";
defparam \Equal4~9 .lut_mask = 64'hFFFFFFFFFFFFFEFF;
defparam \Equal4~9 .shared_arith = "off";

cyclonev_lcell_comb \Equal4~10 (
	.dataa(!\D_iw[0]~q ),
	.datab(!\D_iw[1]~q ),
	.datac(!\D_iw[2]~q ),
	.datad(!\D_iw[3]~q ),
	.datae(!\D_iw[4]~q ),
	.dataf(!\D_iw[5]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal4~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal4~10 .extended_lut = "off";
defparam \Equal4~10 .lut_mask = 64'hFFFFFFFFFFFEFFFF;
defparam \Equal4~10 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_cmp~0 (
	.dataa(!\Equal4~7_combout ),
	.datab(!\Equal4~8_combout ),
	.datac(!\Equal4~9_combout ),
	.datad(!\Equal4~10_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_cmp~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_cmp~0 .extended_lut = "off";
defparam \D_ctrl_cmp~0 .lut_mask = 64'hFFFEFFFEFFFEFFFE;
defparam \D_ctrl_cmp~0 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_cmp~1 (
	.dataa(!\D_iw[12]~q ),
	.datab(!\D_iw[13]~q ),
	.datac(!\Equal4~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_cmp~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_cmp~1 .extended_lut = "off";
defparam \D_ctrl_cmp~1 .lut_mask = 64'hEFEFEFEFEFEFEFEF;
defparam \D_ctrl_cmp~1 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_cmp~2 (
	.dataa(!\D_iw[11]~q ),
	.datab(!\Equal4~5_combout ),
	.datac(!\Equal4~6_combout ),
	.datad(!\D_ctrl_cmp~0_combout ),
	.datae(!\D_ctrl_cmp~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_cmp~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_cmp~2 .extended_lut = "off";
defparam \D_ctrl_cmp~2 .lut_mask = 64'hFFBFFFFFFFBFFFFF;
defparam \D_ctrl_cmp~2 .shared_arith = "off";

dffeas E_ctrl_cmp(
	.clk(clk_clk),
	.d(\D_ctrl_cmp~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_ctrl_cmp~q ),
	.prn(vcc));
defparam E_ctrl_cmp.is_wysiwyg = "true";
defparam E_ctrl_cmp.power_up = "low";

cyclonev_lcell_comb \E_alu_result~0 (
	.dataa(!\E_ctrl_retaddr~q ),
	.datab(!\E_ctrl_logic~q ),
	.datac(!\E_ctrl_cmp~q ),
	.datad(!\E_ctrl_rdctl_inst~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result~0 .extended_lut = "off";
defparam \E_alu_result~0 .lut_mask = 64'hFFFEFFFEFFFEFFFE;
defparam \E_alu_result~0 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_alu_subtract~0 (
	.dataa(!\D_iw[15]~q ),
	.datab(!\D_iw[14]~q ),
	.datac(!\D_iw[11]~q ),
	.datad(!\D_ctrl_cmp~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_alu_subtract~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_alu_subtract~0 .extended_lut = "off";
defparam \D_ctrl_alu_subtract~0 .lut_mask = 64'h96FF96FF96FF96FF;
defparam \D_ctrl_alu_subtract~0 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_alu_subtract~1 (
	.dataa(!\D_iw[4]~q ),
	.datab(!\D_iw[3]~q ),
	.datac(!\D_iw[2]~q ),
	.datad(!\D_iw[1]~q ),
	.datae(!\D_iw[0]~q ),
	.dataf(!\D_ctrl_alu_subtract~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_alu_subtract~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_alu_subtract~1 .extended_lut = "off";
defparam \D_ctrl_alu_subtract~1 .lut_mask = 64'hFFFF6996FFFFFFFF;
defparam \D_ctrl_alu_subtract~1 .shared_arith = "off";

dffeas E_ctrl_alu_subtract(
	.clk(clk_clk),
	.d(\D_ctrl_alu_subtract~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_ctrl_alu_subtract~q ),
	.prn(vcc));
defparam E_ctrl_alu_subtract.is_wysiwyg = "true";
defparam E_ctrl_alu_subtract.power_up = "low";

dffeas \d_readdata_d1[1] (
	.clk(clk_clk),
	.d(d_readdata[1]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d_readdata_d1[1]~q ),
	.prn(vcc));
defparam \d_readdata_d1[1] .is_wysiwyg = "true";
defparam \d_readdata_d1[1] .power_up = "low";

dffeas \d_readdata_d1[17] (
	.clk(clk_clk),
	.d(d_readdata[17]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d_readdata_d1[17]~q ),
	.prn(vcc));
defparam \d_readdata_d1[17] .is_wysiwyg = "true";
defparam \d_readdata_d1[17] .power_up = "low";

dffeas \d_readdata_d1[9] (
	.clk(clk_clk),
	.d(d_readdata[9]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d_readdata_d1[9]~q ),
	.prn(vcc));
defparam \d_readdata_d1[9] .is_wysiwyg = "true";
defparam \d_readdata_d1[9] .power_up = "low";

dffeas \d_readdata_d1[25] (
	.clk(clk_clk),
	.d(d_readdata[25]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d_readdata_d1[25]~q ),
	.prn(vcc));
defparam \d_readdata_d1[25] .is_wysiwyg = "true";
defparam \d_readdata_d1[25] .power_up = "low";

cyclonev_lcell_comb \D_compare_op[1]~0 (
	.dataa(!\D_iw[4]~q ),
	.datab(!\D_iw[15]~q ),
	.datac(!\Equal4~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_compare_op[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_compare_op[1]~0 .extended_lut = "off";
defparam \D_compare_op[1]~0 .lut_mask = 64'h5353535353535353;
defparam \D_compare_op[1]~0 .shared_arith = "off";

dffeas \E_compare_op[1] (
	.clk(clk_clk),
	.d(\D_compare_op[1]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_compare_op[1]~q ),
	.prn(vcc));
defparam \E_compare_op[1] .is_wysiwyg = "true";
defparam \E_compare_op[1] .power_up = "low";

cyclonev_lcell_comb \D_compare_op[0]~1 (
	.dataa(!\D_iw[3]~q ),
	.datab(!\D_iw[14]~q ),
	.datac(!\Equal4~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_compare_op[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_compare_op[0]~1 .extended_lut = "off";
defparam \D_compare_op[0]~1 .lut_mask = 64'h5353535353535353;
defparam \D_compare_op[0]~1 .shared_arith = "off";

dffeas \E_compare_op[0] (
	.clk(clk_clk),
	.d(\D_compare_op[0]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_compare_op[0]~q ),
	.prn(vcc));
defparam \E_compare_op[0] .is_wysiwyg = "true";
defparam \E_compare_op[0] .power_up = "low";

cyclonev_lcell_comb \D_ctrl_a_not_src~0 (
	.dataa(!\D_iw[1]~q ),
	.datab(!\D_iw[2]~q ),
	.datac(!\D_iw[3]~q ),
	.datad(!\D_iw[4]~q ),
	.datae(!\D_iw[5]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_a_not_src~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_a_not_src~0 .extended_lut = "off";
defparam \D_ctrl_a_not_src~0 .lut_mask = 64'hFFFFFFFEFFFFFFFE;
defparam \D_ctrl_a_not_src~0 .shared_arith = "off";

cyclonev_lcell_comb \F_iw[29]~19 (
	.dataa(!\intr_req~0_combout ),
	.datab(!\processor_cpu_ic_data|the_altsyncram|auto_generated|q_b[29] ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[29]~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[29]~19 .extended_lut = "off";
defparam \F_iw[29]~19 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \F_iw[29]~19 .shared_arith = "off";

dffeas \D_iw[29] (
	.clk(clk_clk),
	.d(\F_iw[29]~19_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\F_iw~1_combout ),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\D_iw[29]~q ),
	.prn(vcc));
defparam \D_iw[29] .is_wysiwyg = "true";
defparam \D_iw[29] .power_up = "low";

cyclonev_lcell_comb \F_iw[23]~9 (
	.dataa(!\intr_req~0_combout ),
	.datab(!\processor_cpu_ic_data|the_altsyncram|auto_generated|q_b[23] ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[23]~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[23]~9 .extended_lut = "off";
defparam \F_iw[23]~9 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \F_iw[23]~9 .shared_arith = "off";

dffeas \D_iw[23] (
	.clk(clk_clk),
	.d(\F_iw[23]~9_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\F_iw~1_combout ),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\D_iw[23]~q ),
	.prn(vcc));
defparam \D_iw[23] .is_wysiwyg = "true";
defparam \D_iw[23] .power_up = "low";

cyclonev_lcell_comb \F_iw[18]~30 (
	.dataa(!\F_iw~1_combout ),
	.datab(!\intr_req~0_combout ),
	.datac(!\processor_cpu_ic_data|the_altsyncram|auto_generated|q_b[18] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[18]~30_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[18]~30 .extended_lut = "off";
defparam \F_iw[18]~30 .lut_mask = 64'hDFDFDFDFDFDFDFDF;
defparam \F_iw[18]~30 .shared_arith = "off";

dffeas \D_iw[18] (
	.clk(clk_clk),
	.d(\F_iw[18]~30_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\D_iw[18]~q ),
	.prn(vcc));
defparam \D_iw[18] .is_wysiwyg = "true";
defparam \D_iw[18] .power_up = "low";

cyclonev_lcell_comb \D_ctrl_implicit_dst_eretaddr~1 (
	.dataa(!\D_iw[11]~q ),
	.datab(!\D_iw[12]~q ),
	.datac(!\D_iw[13]~q ),
	.datad(!\D_iw[14]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_implicit_dst_eretaddr~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_implicit_dst_eretaddr~1 .extended_lut = "off";
defparam \D_ctrl_implicit_dst_eretaddr~1 .lut_mask = 64'hFFDFFFDFFFDFFFDF;
defparam \D_ctrl_implicit_dst_eretaddr~1 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_implicit_dst_eretaddr~2 (
	.dataa(!\D_iw[16]~q ),
	.datab(!\D_iw[15]~q ),
	.datac(!\Equal4~0_combout ),
	.datad(!\D_ctrl_implicit_dst_eretaddr~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_implicit_dst_eretaddr~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_implicit_dst_eretaddr~2 .extended_lut = "off";
defparam \D_ctrl_implicit_dst_eretaddr~2 .lut_mask = 64'hDFFFDFFFDFFFDFFF;
defparam \D_ctrl_implicit_dst_eretaddr~2 .shared_arith = "off";

cyclonev_lcell_comb \D_dst_regnum[1]~2 (
	.dataa(!\D_iw[23]~q ),
	.datab(!\D_ctrl_b_not_src~0_combout ),
	.datac(!\D_ctrl_implicit_dst_retaddr~0_combout ),
	.datad(!\D_iw[18]~q ),
	.datae(!\D_ctrl_implicit_dst_eretaddr~2_combout ),
	.dataf(!\D_ctrl_implicit_dst_eretaddr~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_dst_regnum[1]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_dst_regnum[1]~2 .extended_lut = "off";
defparam \D_dst_regnum[1]~2 .lut_mask = 64'hDFFF1FFFFFFFFFFF;
defparam \D_dst_regnum[1]~2 .shared_arith = "off";

cyclonev_lcell_comb \F_iw[22]~8 (
	.dataa(!\processor_cpu_ic_data|the_altsyncram|auto_generated|q_b[22] ),
	.datab(!\intr_req~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[22]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[22]~8 .extended_lut = "off";
defparam \F_iw[22]~8 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \F_iw[22]~8 .shared_arith = "off";

dffeas \D_iw[22] (
	.clk(clk_clk),
	.d(\F_iw[22]~8_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\F_iw~1_combout ),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\D_iw[22]~q ),
	.prn(vcc));
defparam \D_iw[22] .is_wysiwyg = "true";
defparam \D_iw[22] .power_up = "low";

cyclonev_lcell_comb \F_iw[17]~31 (
	.dataa(!\intr_req~0_combout ),
	.datab(!\processor_cpu_ic_data|the_altsyncram|auto_generated|q_b[17] ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[17]~31_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[17]~31 .extended_lut = "off";
defparam \F_iw[17]~31 .lut_mask = 64'h7777777777777777;
defparam \F_iw[17]~31 .shared_arith = "off";

dffeas \D_iw[17] (
	.clk(clk_clk),
	.d(\F_iw[17]~31_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\F_iw~1_combout ),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\D_iw[17]~q ),
	.prn(vcc));
defparam \D_iw[17] .is_wysiwyg = "true";
defparam \D_iw[17] .power_up = "low";

cyclonev_lcell_comb \D_dst_regnum[4]~0 (
	.dataa(!\D_ctrl_implicit_dst_retaddr~0_combout ),
	.datab(!\D_iw[15]~q ),
	.datac(!\D_iw[14]~q ),
	.datad(!\Equal4~1_combout ),
	.datae(!\Equal107~0_combout ),
	.dataf(!\D_ctrl_implicit_dst_eretaddr~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_dst_regnum[4]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_dst_regnum[4]~0 .extended_lut = "off";
defparam \D_dst_regnum[4]~0 .lut_mask = 64'hFFFFFFFFFFFFFFEF;
defparam \D_dst_regnum[4]~0 .shared_arith = "off";

cyclonev_lcell_comb \D_dst_regnum[0]~3 (
	.dataa(!\D_iw[22]~q ),
	.datab(!\D_ctrl_b_not_src~0_combout ),
	.datac(!\D_iw[17]~q ),
	.datad(!\D_dst_regnum[4]~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_dst_regnum[0]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_dst_regnum[0]~3 .extended_lut = "off";
defparam \D_dst_regnum[0]~3 .lut_mask = 64'hDF1FDF1FDF1FDF1F;
defparam \D_dst_regnum[0]~3 .shared_arith = "off";

cyclonev_lcell_comb \F_iw[25]~10 (
	.dataa(!\intr_req~0_combout ),
	.datab(!\processor_cpu_ic_data|the_altsyncram|auto_generated|q_b[25] ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[25]~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[25]~10 .extended_lut = "off";
defparam \F_iw[25]~10 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \F_iw[25]~10 .shared_arith = "off";

dffeas \D_iw[25] (
	.clk(clk_clk),
	.d(\F_iw[25]~10_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\F_iw~1_combout ),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\D_iw[25]~q ),
	.prn(vcc));
defparam \D_iw[25] .is_wysiwyg = "true";
defparam \D_iw[25] .power_up = "low";

cyclonev_lcell_comb \F_iw[20]~28 (
	.dataa(!\F_iw~1_combout ),
	.datab(!\intr_req~0_combout ),
	.datac(!\processor_cpu_ic_data|the_altsyncram|auto_generated|q_b[20] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[20]~28_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[20]~28 .extended_lut = "off";
defparam \F_iw[20]~28 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \F_iw[20]~28 .shared_arith = "off";

dffeas \D_iw[20] (
	.clk(clk_clk),
	.d(\F_iw[20]~28_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\D_iw[20]~q ),
	.prn(vcc));
defparam \D_iw[20] .is_wysiwyg = "true";
defparam \D_iw[20] .power_up = "low";

cyclonev_lcell_comb \D_dst_regnum[3]~4 (
	.dataa(!\D_iw[25]~q ),
	.datab(!\D_ctrl_b_not_src~0_combout ),
	.datac(!\D_iw[20]~q ),
	.datad(!\D_dst_regnum[4]~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_dst_regnum[3]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_dst_regnum[3]~4 .extended_lut = "off";
defparam \D_dst_regnum[3]~4 .lut_mask = 64'hDF1FDF1FDF1FDF1F;
defparam \D_dst_regnum[3]~4 .shared_arith = "off";

cyclonev_lcell_comb \F_iw[26]~11 (
	.dataa(!\intr_req~0_combout ),
	.datab(!\processor_cpu_ic_data|the_altsyncram|auto_generated|q_b[26] ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[26]~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[26]~11 .extended_lut = "off";
defparam \F_iw[26]~11 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \F_iw[26]~11 .shared_arith = "off";

dffeas \D_iw[26] (
	.clk(clk_clk),
	.d(\F_iw[26]~11_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\F_iw~1_combout ),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\D_iw[26]~q ),
	.prn(vcc));
defparam \D_iw[26] .is_wysiwyg = "true";
defparam \D_iw[26] .power_up = "low";

cyclonev_lcell_comb \F_iw[21]~18 (
	.dataa(!\F_iw~1_combout ),
	.datab(!\intr_req~0_combout ),
	.datac(!\processor_cpu_ic_data|the_altsyncram|auto_generated|q_b[21] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[21]~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[21]~18 .extended_lut = "off";
defparam \F_iw[21]~18 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \F_iw[21]~18 .shared_arith = "off";

dffeas \D_iw[21] (
	.clk(clk_clk),
	.d(\F_iw[21]~18_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\D_iw[21]~q ),
	.prn(vcc));
defparam \D_iw[21] .is_wysiwyg = "true";
defparam \D_iw[21] .power_up = "low";

cyclonev_lcell_comb \D_dst_regnum[4]~5 (
	.dataa(!\D_iw[26]~q ),
	.datab(!\D_ctrl_b_not_src~0_combout ),
	.datac(!\D_iw[21]~q ),
	.datad(!\D_dst_regnum[4]~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_dst_regnum[4]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_dst_regnum[4]~5 .extended_lut = "off";
defparam \D_dst_regnum[4]~5 .lut_mask = 64'hDF1FDF1FDF1FDF1F;
defparam \D_dst_regnum[4]~5 .shared_arith = "off";

cyclonev_lcell_comb \D_wr_dst_reg~0 (
	.dataa(!\D_valid~combout ),
	.datab(!\D_iw[2]~q ),
	.datac(!\D_iw[1]~q ),
	.datad(!\D_iw[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_wr_dst_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_wr_dst_reg~0 .extended_lut = "off";
defparam \D_wr_dst_reg~0 .lut_mask = 64'hDFFDDFFDDFFDDFFD;
defparam \D_wr_dst_reg~0 .shared_arith = "off";

cyclonev_lcell_comb D_wr_dst_reg(
	.dataa(!\D_dst_regnum[1]~2_combout ),
	.datab(!\D_dst_regnum[0]~3_combout ),
	.datac(!\D_dst_regnum[2]~1_combout ),
	.datad(!\D_dst_regnum[3]~4_combout ),
	.datae(!\D_dst_regnum[4]~5_combout ),
	.dataf(!\D_wr_dst_reg~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_wr_dst_reg~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam D_wr_dst_reg.extended_lut = "off";
defparam D_wr_dst_reg.lut_mask = 64'h7FFFFFFFFFFFFFFF;
defparam D_wr_dst_reg.shared_arith = "off";

dffeas E_wr_dst_reg_from_D(
	.clk(clk_clk),
	.d(\D_wr_dst_reg~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_wr_dst_reg_from_D~q ),
	.prn(vcc));
defparam E_wr_dst_reg_from_D.is_wysiwyg = "true";
defparam E_wr_dst_reg_from_D.power_up = "low";

cyclonev_lcell_comb \E_wr_dst_reg~0 (
	.dataa(!\M_pipe_flush~q ),
	.datab(!\E_hbreak_req~combout ),
	.datac(!\E_wr_dst_reg_from_D~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_wr_dst_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_wr_dst_reg~0 .extended_lut = "off";
defparam \E_wr_dst_reg~0 .lut_mask = 64'hFBFBFBFBFBFBFBFB;
defparam \E_wr_dst_reg~0 .shared_arith = "off";

dffeas \E_dst_regnum[0] (
	.clk(clk_clk),
	.d(\D_dst_regnum[0]~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_dst_regnum[0]~q ),
	.prn(vcc));
defparam \E_dst_regnum[0] .is_wysiwyg = "true";
defparam \E_dst_regnum[0] .power_up = "low";

dffeas \E_dst_regnum[1] (
	.clk(clk_clk),
	.d(\D_dst_regnum[1]~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_dst_regnum[1]~q ),
	.prn(vcc));
defparam \E_dst_regnum[1] .is_wysiwyg = "true";
defparam \E_dst_regnum[1] .power_up = "low";

cyclonev_lcell_comb \F_iw[27]~20 (
	.dataa(!\intr_req~0_combout ),
	.datab(!\processor_cpu_ic_data|the_altsyncram|auto_generated|q_b[27] ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[27]~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[27]~20 .extended_lut = "off";
defparam \F_iw[27]~20 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \F_iw[27]~20 .shared_arith = "off";

dffeas \D_iw[27] (
	.clk(clk_clk),
	.d(\F_iw[27]~20_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\F_iw~1_combout ),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\D_iw[27]~q ),
	.prn(vcc));
defparam \D_iw[27] .is_wysiwyg = "true";
defparam \D_iw[27] .power_up = "low";

cyclonev_lcell_comb \F_iw[28]~21 (
	.dataa(!\intr_req~0_combout ),
	.datab(!\processor_cpu_ic_data|the_altsyncram|auto_generated|q_b[28] ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[28]~21_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[28]~21 .extended_lut = "off";
defparam \F_iw[28]~21 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \F_iw[28]~21 .shared_arith = "off";

dffeas \D_iw[28] (
	.clk(clk_clk),
	.d(\F_iw[28]~21_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\F_iw~1_combout ),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\D_iw[28]~q ),
	.prn(vcc));
defparam \D_iw[28] .is_wysiwyg = "true";
defparam \D_iw[28] .power_up = "low";

cyclonev_lcell_comb \D_src1_hazard_E~0 (
	.dataa(!\E_dst_regnum[0]~q ),
	.datab(!\E_dst_regnum[1]~q ),
	.datac(!\D_iw[27]~q ),
	.datad(!\D_iw[28]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_hazard_E~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src1_hazard_E~0 .extended_lut = "off";
defparam \D_src1_hazard_E~0 .lut_mask = 64'h6996699669966996;
defparam \D_src1_hazard_E~0 .shared_arith = "off";

dffeas \E_dst_regnum[3] (
	.clk(clk_clk),
	.d(\D_dst_regnum[3]~4_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_dst_regnum[3]~q ),
	.prn(vcc));
defparam \E_dst_regnum[3] .is_wysiwyg = "true";
defparam \E_dst_regnum[3] .power_up = "low";

dffeas \E_dst_regnum[4] (
	.clk(clk_clk),
	.d(\D_dst_regnum[4]~5_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_dst_regnum[4]~q ),
	.prn(vcc));
defparam \E_dst_regnum[4] .is_wysiwyg = "true";
defparam \E_dst_regnum[4] .power_up = "low";

cyclonev_lcell_comb \F_iw[30]~22 (
	.dataa(!\intr_req~0_combout ),
	.datab(!\processor_cpu_ic_data|the_altsyncram|auto_generated|q_b[30] ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[30]~22_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[30]~22 .extended_lut = "off";
defparam \F_iw[30]~22 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \F_iw[30]~22 .shared_arith = "off";

dffeas \D_iw[30] (
	.clk(clk_clk),
	.d(\F_iw[30]~22_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\F_iw~1_combout ),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\D_iw[30]~q ),
	.prn(vcc));
defparam \D_iw[30] .is_wysiwyg = "true";
defparam \D_iw[30] .power_up = "low";

cyclonev_lcell_comb \F_iw[31]~23 (
	.dataa(!\intr_req~0_combout ),
	.datab(!\processor_cpu_ic_data|the_altsyncram|auto_generated|q_b[31] ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[31]~23_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[31]~23 .extended_lut = "off";
defparam \F_iw[31]~23 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \F_iw[31]~23 .shared_arith = "off";

dffeas \D_iw[31] (
	.clk(clk_clk),
	.d(\F_iw[31]~23_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\F_iw~1_combout ),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\D_iw[31]~q ),
	.prn(vcc));
defparam \D_iw[31] .is_wysiwyg = "true";
defparam \D_iw[31] .power_up = "low";

cyclonev_lcell_comb \D_src1_hazard_E~1 (
	.dataa(!\E_dst_regnum[3]~q ),
	.datab(!\E_dst_regnum[4]~q ),
	.datac(!\D_iw[30]~q ),
	.datad(!\D_iw[31]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_hazard_E~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src1_hazard_E~1 .extended_lut = "off";
defparam \D_src1_hazard_E~1 .lut_mask = 64'h6996699669966996;
defparam \D_src1_hazard_E~1 .shared_arith = "off";

cyclonev_lcell_comb D_src1_hazard_E(
	.dataa(!\E_dst_regnum[2]~q ),
	.datab(!\D_ctrl_a_not_src~0_combout ),
	.datac(!\D_iw[29]~q ),
	.datad(!\E_wr_dst_reg~0_combout ),
	.datae(!\D_src1_hazard_E~0_combout ),
	.dataf(!\D_src1_hazard_E~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_hazard_E~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam D_src1_hazard_E.extended_lut = "off";
defparam D_src1_hazard_E.lut_mask = 64'hFFDEFFFFFFFFFFFF;
defparam D_src1_hazard_E.shared_arith = "off";

dffeas E_src1_hazard_M(
	.clk(clk_clk),
	.d(\D_src1_hazard_E~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_src1_hazard_M~q ),
	.prn(vcc));
defparam E_src1_hazard_M.is_wysiwyg = "true";
defparam E_src1_hazard_M.power_up = "low";

cyclonev_lcell_comb \D_ctrl_shift_rot_right~0 (
	.dataa(!\D_iw[14]~q ),
	.datab(!\D_ctrl_shift_logical~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_shift_rot_right~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_shift_rot_right~0 .extended_lut = "off";
defparam \D_ctrl_shift_rot_right~0 .lut_mask = 64'h7777777777777777;
defparam \D_ctrl_shift_rot_right~0 .shared_arith = "off";

dffeas E_ctrl_shift_rot_right(
	.clk(clk_clk),
	.d(\D_ctrl_shift_rot_right~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_ctrl_shift_rot_right~q ),
	.prn(vcc));
defparam E_ctrl_shift_rot_right.is_wysiwyg = "true";
defparam E_ctrl_shift_rot_right.power_up = "low";

dffeas M_ctrl_shift_rot_right(
	.clk(clk_clk),
	.d(\E_ctrl_shift_rot_right~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\M_ctrl_shift_rot_right~q ),
	.prn(vcc));
defparam M_ctrl_shift_rot_right.is_wysiwyg = "true";
defparam M_ctrl_shift_rot_right.power_up = "low";

cyclonev_lcell_comb \D_ctrl_shift_logical~1 (
	.dataa(!\D_iw[16]~q ),
	.datab(!\D_iw[15]~q ),
	.datac(!\D_ctrl_shift_logical~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_shift_logical~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_shift_logical~1 .extended_lut = "off";
defparam \D_ctrl_shift_logical~1 .lut_mask = 64'hBFBFBFBFBFBFBFBF;
defparam \D_ctrl_shift_logical~1 .shared_arith = "off";

dffeas E_ctrl_shift_logical(
	.clk(clk_clk),
	.d(\D_ctrl_shift_logical~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_ctrl_shift_logical~q ),
	.prn(vcc));
defparam E_ctrl_shift_logical.is_wysiwyg = "true";
defparam E_ctrl_shift_logical.power_up = "low";

dffeas M_ctrl_shift_logical(
	.clk(clk_clk),
	.d(\E_ctrl_shift_logical~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\M_ctrl_shift_logical~q ),
	.prn(vcc));
defparam M_ctrl_shift_logical.is_wysiwyg = "true";
defparam M_ctrl_shift_logical.power_up = "low";

cyclonev_lcell_comb \D_ctrl_rot_right~0 (
	.dataa(!\D_iw[15]~q ),
	.datab(!\D_iw[14]~q ),
	.datac(!\D_ctrl_shift_logical~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_rot_right~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_rot_right~0 .extended_lut = "off";
defparam \D_ctrl_rot_right~0 .lut_mask = 64'hBFBFBFBFBFBFBFBF;
defparam \D_ctrl_rot_right~0 .shared_arith = "off";

dffeas E_ctrl_rot_right(
	.clk(clk_clk),
	.d(\D_ctrl_rot_right~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_ctrl_rot_right~q ),
	.prn(vcc));
defparam E_ctrl_rot_right.is_wysiwyg = "true";
defparam E_ctrl_rot_right.power_up = "low";

dffeas M_ctrl_rot_right(
	.clk(clk_clk),
	.d(\E_ctrl_rot_right~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\M_ctrl_rot_right~q ),
	.prn(vcc));
defparam M_ctrl_rot_right.is_wysiwyg = "true";
defparam M_ctrl_rot_right.power_up = "low";

cyclonev_lcell_comb \M_shift_rot_fill_bit~0 (
	.dataa(!\M_shift_rot_result[0]~q ),
	.datab(!\M_ctrl_shift_logical~q ),
	.datac(!\M_ctrl_rot_right~q ),
	.datad(!\M_shift_rot_result[31]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_shift_rot_fill_bit~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_shift_rot_fill_bit~0 .extended_lut = "off";
defparam \M_shift_rot_fill_bit~0 .lut_mask = 64'hC5FFC5FFC5FFC5FF;
defparam \M_shift_rot_fill_bit~0 .shared_arith = "off";

dffeas \d_readdata_d1[31] (
	.clk(clk_clk),
	.d(d_readdata[31]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d_readdata_d1[31]~q ),
	.prn(vcc));
defparam \d_readdata_d1[31] .is_wysiwyg = "true";
defparam \d_readdata_d1[31] .power_up = "low";

dffeas \d_readdata_d1[15] (
	.clk(clk_clk),
	.d(d_readdata[15]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d_readdata_d1[15]~q ),
	.prn(vcc));
defparam \d_readdata_d1[15] .is_wysiwyg = "true";
defparam \d_readdata_d1[15] .power_up = "low";

dffeas \d_readdata_d1[23] (
	.clk(clk_clk),
	.d(d_readdata[23]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d_readdata_d1[23]~q ),
	.prn(vcc));
defparam \d_readdata_d1[23] .is_wysiwyg = "true";
defparam \d_readdata_d1[23] .power_up = "low";

dffeas \M_iw[4] (
	.clk(clk_clk),
	.d(\E_iw[4]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\M_iw[4]~q ),
	.prn(vcc));
defparam \M_iw[4] .is_wysiwyg = "true";
defparam \M_iw[4] .power_up = "low";

dffeas \M_iw[3] (
	.clk(clk_clk),
	.d(\E_iw[3]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\M_iw[3]~q ),
	.prn(vcc));
defparam \M_iw[3] .is_wysiwyg = "true";
defparam \M_iw[3] .power_up = "low";

cyclonev_lcell_comb \av_sign_bit~0 (
	.dataa(!\M_alu_result[0]~q ),
	.datab(!\M_iw[4]~q ),
	.datac(!\M_iw[3]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_sign_bit~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_sign_bit~0 .extended_lut = "off";
defparam \av_sign_bit~0 .lut_mask = 64'hDFDFDFDFDFDFDFDF;
defparam \av_sign_bit~0 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_b_is_dst~0 (
	.dataa(!\D_iw[0]~q ),
	.datab(!\D_iw[1]~q ),
	.datac(!\D_iw[2]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_b_is_dst~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_b_is_dst~0 .extended_lut = "off";
defparam \D_ctrl_b_is_dst~0 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \D_ctrl_b_is_dst~0 .shared_arith = "off";

dffeas E_ctrl_ld_signed(
	.clk(clk_clk),
	.d(\D_ctrl_b_is_dst~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_ctrl_ld_signed~q ),
	.prn(vcc));
defparam E_ctrl_ld_signed.is_wysiwyg = "true";
defparam E_ctrl_ld_signed.power_up = "low";

dffeas M_ctrl_ld_signed(
	.clk(clk_clk),
	.d(\E_ctrl_ld_signed~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\M_ctrl_ld_signed~q ),
	.prn(vcc));
defparam M_ctrl_ld_signed.is_wysiwyg = "true";
defparam M_ctrl_ld_signed.power_up = "low";

dffeas \d_readdata_d1[7] (
	.clk(clk_clk),
	.d(d_readdata[7]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d_readdata_d1[7]~q ),
	.prn(vcc));
defparam \d_readdata_d1[7] .is_wysiwyg = "true";
defparam \d_readdata_d1[7] .power_up = "low";

cyclonev_lcell_comb \av_fill_bit~0 (
	.dataa(!\M_alu_result[1]~q ),
	.datab(!\d_readdata_d1[31]~q ),
	.datac(!\d_readdata_d1[15]~q ),
	.datad(!\d_readdata_d1[23]~q ),
	.datae(!\av_sign_bit~0_combout ),
	.dataf(!\M_ctrl_ld_signed~q ),
	.datag(!\d_readdata_d1[7]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_fill_bit~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_fill_bit~0 .extended_lut = "on";
defparam \av_fill_bit~0 .lut_mask = 64'hFFD8FFD8FFD8FFD8;
defparam \av_fill_bit~0 .shared_arith = "off";

dffeas \d_readdata_d1[30] (
	.clk(clk_clk),
	.d(d_readdata[30]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d_readdata_d1[30]~q ),
	.prn(vcc));
defparam \d_readdata_d1[30] .is_wysiwyg = "true";
defparam \d_readdata_d1[30] .power_up = "low";

dffeas \av_ld_data_aligned_or_div[30] (
	.clk(clk_clk),
	.d(\av_fill_bit~0_combout ),
	.asdata(\d_readdata_d1[30]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\M_iw[4]~q ),
	.ena(vcc),
	.q(\av_ld_data_aligned_or_div[30]~q ),
	.prn(vcc));
defparam \av_ld_data_aligned_or_div[30] .is_wysiwyg = "true";
defparam \av_ld_data_aligned_or_div[30] .power_up = "low";

cyclonev_lcell_comb \E_stw_data[30]~15 (
	.dataa(!\E_src2_hazard_M~q ),
	.datab(!\M_ctrl_shift_rot~q ),
	.datac(!\av_ld_or_div_done~q ),
	.datad(!\M_shift_rot_result[30]~q ),
	.datae(!\av_ld_data_aligned_or_div[30]~q ),
	.dataf(!\M_alu_result[30]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_stw_data[30]~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_stw_data[30]~15 .extended_lut = "off";
defparam \E_stw_data[30]~15 .lut_mask = 64'h7DFFFFFFFFFFFFFF;
defparam \E_stw_data[30]~15 .shared_arith = "off";

cyclonev_lcell_comb \M_wr_data_unfiltered[30]~19 (
	.dataa(!\M_ctrl_shift_rot~q ),
	.datab(!\av_ld_or_div_done~q ),
	.datac(!\M_shift_rot_result[30]~q ),
	.datad(!\av_ld_data_aligned_or_div[30]~q ),
	.datae(!\M_alu_result[30]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_wr_data_unfiltered[30]~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_wr_data_unfiltered[30]~19 .extended_lut = "off";
defparam \M_wr_data_unfiltered[30]~19 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \M_wr_data_unfiltered[30]~19 .shared_arith = "off";

dffeas \M_dst_regnum[4] (
	.clk(clk_clk),
	.d(\E_dst_regnum[4]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\M_dst_regnum[4]~q ),
	.prn(vcc));
defparam \M_dst_regnum[4] .is_wysiwyg = "true";
defparam \M_dst_regnum[4] .power_up = "low";

dffeas M_wr_dst_reg(
	.clk(clk_clk),
	.d(\E_wr_dst_reg~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\M_wr_dst_reg~q ),
	.prn(vcc));
defparam M_wr_dst_reg.is_wysiwyg = "true";
defparam M_wr_dst_reg.power_up = "low";

dffeas \M_dst_regnum[0] (
	.clk(clk_clk),
	.d(\E_dst_regnum[0]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\M_dst_regnum[0]~q ),
	.prn(vcc));
defparam \M_dst_regnum[0] .is_wysiwyg = "true";
defparam \M_dst_regnum[0] .power_up = "low";

dffeas \M_dst_regnum[1] (
	.clk(clk_clk),
	.d(\E_dst_regnum[1]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\M_dst_regnum[1]~q ),
	.prn(vcc));
defparam \M_dst_regnum[1] .is_wysiwyg = "true";
defparam \M_dst_regnum[1] .power_up = "low";

cyclonev_lcell_comb \D_src2_hazard_M~0 (
	.dataa(!\D_iw[22]~q ),
	.datab(!\D_iw[23]~q ),
	.datac(!\M_wr_dst_reg~q ),
	.datad(!\M_dst_regnum[0]~q ),
	.datae(!\M_dst_regnum[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_hazard_M~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_hazard_M~0 .extended_lut = "off";
defparam \D_src2_hazard_M~0 .lut_mask = 64'hF6F9F9F6F6F9F9F6;
defparam \D_src2_hazard_M~0 .shared_arith = "off";

dffeas \M_dst_regnum[2] (
	.clk(clk_clk),
	.d(\E_dst_regnum[2]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\M_dst_regnum[2]~q ),
	.prn(vcc));
defparam \M_dst_regnum[2] .is_wysiwyg = "true";
defparam \M_dst_regnum[2] .power_up = "low";

dffeas \M_dst_regnum[3] (
	.clk(clk_clk),
	.d(\E_dst_regnum[3]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\M_dst_regnum[3]~q ),
	.prn(vcc));
defparam \M_dst_regnum[3] .is_wysiwyg = "true";
defparam \M_dst_regnum[3] .power_up = "low";

cyclonev_lcell_comb \D_src2_hazard_M~1 (
	.dataa(!\D_iw[24]~q ),
	.datab(!\D_iw[25]~q ),
	.datac(!\M_dst_regnum[2]~q ),
	.datad(!\M_dst_regnum[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_hazard_M~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_hazard_M~1 .extended_lut = "off";
defparam \D_src2_hazard_M~1 .lut_mask = 64'h6996699669966996;
defparam \D_src2_hazard_M~1 .shared_arith = "off";

cyclonev_lcell_comb D_src2_hazard_M(
	.dataa(!\D_iw[26]~q ),
	.datab(!\M_dst_regnum[4]~q ),
	.datac(!\D_ctrl_b_not_src~0_combout ),
	.datad(!\D_src2_hazard_M~0_combout ),
	.datae(!\D_src2_hazard_M~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_hazard_M~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam D_src2_hazard_M.extended_lut = "off";
defparam D_src2_hazard_M.lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam D_src2_hazard_M.shared_arith = "off";

dffeas \W_dst_regnum[4] (
	.clk(clk_clk),
	.d(\M_dst_regnum[4]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\W_dst_regnum[4]~q ),
	.prn(vcc));
defparam \W_dst_regnum[4] .is_wysiwyg = "true";
defparam \W_dst_regnum[4] .power_up = "low";

cyclonev_lcell_comb \W_wr_dst_reg~0 (
	.dataa(!\M_wr_dst_reg~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\W_wr_dst_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \W_wr_dst_reg~0 .extended_lut = "off";
defparam \W_wr_dst_reg~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \W_wr_dst_reg~0 .shared_arith = "off";

dffeas W_wr_dst_reg(
	.clk(clk_clk),
	.d(\W_wr_dst_reg~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\W_wr_dst_reg~q ),
	.prn(vcc));
defparam W_wr_dst_reg.is_wysiwyg = "true";
defparam W_wr_dst_reg.power_up = "low";

dffeas \W_dst_regnum[0] (
	.clk(clk_clk),
	.d(\M_dst_regnum[0]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\W_dst_regnum[0]~q ),
	.prn(vcc));
defparam \W_dst_regnum[0] .is_wysiwyg = "true";
defparam \W_dst_regnum[0] .power_up = "low";

dffeas \W_dst_regnum[1] (
	.clk(clk_clk),
	.d(\M_dst_regnum[1]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\W_dst_regnum[1]~q ),
	.prn(vcc));
defparam \W_dst_regnum[1] .is_wysiwyg = "true";
defparam \W_dst_regnum[1] .power_up = "low";

cyclonev_lcell_comb \D_src2_hazard_W~0 (
	.dataa(!\D_iw[22]~q ),
	.datab(!\D_iw[23]~q ),
	.datac(!\W_wr_dst_reg~q ),
	.datad(!\W_dst_regnum[0]~q ),
	.datae(!\W_dst_regnum[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_hazard_W~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_hazard_W~0 .extended_lut = "off";
defparam \D_src2_hazard_W~0 .lut_mask = 64'h6F9F9F6F6F9F9F6F;
defparam \D_src2_hazard_W~0 .shared_arith = "off";

dffeas \W_dst_regnum[2] (
	.clk(clk_clk),
	.d(\M_dst_regnum[2]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\W_dst_regnum[2]~q ),
	.prn(vcc));
defparam \W_dst_regnum[2] .is_wysiwyg = "true";
defparam \W_dst_regnum[2] .power_up = "low";

dffeas \W_dst_regnum[3] (
	.clk(clk_clk),
	.d(\M_dst_regnum[3]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\W_dst_regnum[3]~q ),
	.prn(vcc));
defparam \W_dst_regnum[3] .is_wysiwyg = "true";
defparam \W_dst_regnum[3] .power_up = "low";

cyclonev_lcell_comb \D_src2_hazard_W~1 (
	.dataa(!\D_iw[24]~q ),
	.datab(!\D_iw[25]~q ),
	.datac(!\W_dst_regnum[2]~q ),
	.datad(!\W_dst_regnum[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_hazard_W~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_hazard_W~1 .extended_lut = "off";
defparam \D_src2_hazard_W~1 .lut_mask = 64'h6996699669966996;
defparam \D_src2_hazard_W~1 .shared_arith = "off";

cyclonev_lcell_comb D_src2_hazard_W(
	.dataa(!\D_iw[26]~q ),
	.datab(!\D_ctrl_b_not_src~0_combout ),
	.datac(!\W_dst_regnum[4]~q ),
	.datad(!\D_src2_hazard_W~0_combout ),
	.datae(!\D_src2_hazard_W~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_hazard_W~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam D_src2_hazard_W.extended_lut = "off";
defparam D_src2_hazard_W.lut_mask = 64'h7BFFFFFF7BFFFFFF;
defparam D_src2_hazard_W.shared_arith = "off";

dffeas \W_wr_data[30] (
	.clk(clk_clk),
	.d(\M_wr_data_unfiltered[30]~19_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\W_wr_data[30]~q ),
	.prn(vcc));
defparam \W_wr_data[30] .is_wysiwyg = "true";
defparam \W_wr_data[30] .power_up = "low";

cyclonev_lcell_comb \D_src2_prelim[30]~19 (
	.dataa(!\M_wr_data_unfiltered[30]~19_combout ),
	.datab(!\D_src2_hazard_M~combout ),
	.datac(!\D_src2_hazard_W~combout ),
	.datad(!\W_wr_data[30]~q ),
	.datae(!\processor_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[30] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_prelim[30]~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_prelim[30]~19 .extended_lut = "off";
defparam \D_src2_prelim[30]~19 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \D_src2_prelim[30]~19 .shared_arith = "off";

dffeas \E_src2_prelim[30] (
	.clk(clk_clk),
	.d(\D_src2_prelim[30]~19_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_src2_prelim[30]~q ),
	.prn(vcc));
defparam \E_src2_prelim[30] .is_wysiwyg = "true";
defparam \E_src2_prelim[30] .power_up = "low";

cyclonev_lcell_comb \E_stw_data[30]~16 (
	.dataa(!\E_src2_hazard_M~q ),
	.datab(!\E_src2_prelim[30]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_stw_data[30]~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_stw_data[30]~16 .extended_lut = "off";
defparam \E_stw_data[30]~16 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \E_stw_data[30]~16 .shared_arith = "off";

cyclonev_lcell_comb \E_stw_data[30]~17 (
	.dataa(!\E_stw_data[30]~15_combout ),
	.datab(!\E_stw_data[30]~16_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_stw_data[30]~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_stw_data[30]~17 .extended_lut = "off";
defparam \E_stw_data[30]~17 .lut_mask = 64'h7777777777777777;
defparam \E_stw_data[30]~17 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_logic~1 (
	.dataa(!\D_iw[5]~q ),
	.datab(!\D_iw[4]~q ),
	.datac(!\D_iw[3]~q ),
	.datad(!\D_iw[2]~q ),
	.datae(!\D_iw[1]~q ),
	.dataf(!\D_iw[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_logic~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_logic~1 .extended_lut = "off";
defparam \D_ctrl_logic~1 .lut_mask = 64'hFFFFFFFFFFFFBFFF;
defparam \D_ctrl_logic~1 .shared_arith = "off";

cyclonev_lcell_comb D_ctrl_unsigned_lo_imm16(
	.dataa(!\D_iw[11]~q ),
	.datab(!\Equal4~7_combout ),
	.datac(!\Equal4~8_combout ),
	.datad(!\D_ctrl_shift_logical~0_combout ),
	.datae(!\D_ctrl_logic~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_unsigned_lo_imm16~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam D_ctrl_unsigned_lo_imm16.extended_lut = "off";
defparam D_ctrl_unsigned_lo_imm16.lut_mask = 64'hBFFFFFFFBFFFFFFF;
defparam D_ctrl_unsigned_lo_imm16.shared_arith = "off";

cyclonev_lcell_comb \Equal171~0 (
	.dataa(!\D_iw[11]~q ),
	.datab(!\Equal4~7_combout ),
	.datac(!\Equal4~8_combout ),
	.datad(!\D_ctrl_shift_logical~0_combout ),
	.datae(!\D_ctrl_hi_imm16~0_combout ),
	.dataf(!\D_ctrl_logic~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal171~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal171~0 .extended_lut = "off";
defparam \Equal171~0 .lut_mask = 64'hBFFFFFFFFFFFFFFF;
defparam \Equal171~0 .shared_arith = "off";

dffeas \E_src2_imm[30] (
	.clk(clk_clk),
	.d(\D_iw[21]~q ),
	.asdata(\D_iw[20]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\D_ctrl_unsigned_lo_imm16~combout ),
	.sload(\Equal171~0_combout ),
	.ena(\W_stall~combout ),
	.q(\E_src2_imm[30]~q ),
	.prn(vcc));
defparam \E_src2_imm[30] .is_wysiwyg = "true";
defparam \E_src2_imm[30] .power_up = "low";

dffeas \d_readdata_d1[28] (
	.clk(clk_clk),
	.d(d_readdata[28]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d_readdata_d1[28]~q ),
	.prn(vcc));
defparam \d_readdata_d1[28] .is_wysiwyg = "true";
defparam \d_readdata_d1[28] .power_up = "low";

dffeas \av_ld_data_aligned_or_div[28] (
	.clk(clk_clk),
	.d(\av_fill_bit~0_combout ),
	.asdata(\d_readdata_d1[28]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\M_iw[4]~q ),
	.ena(vcc),
	.q(\av_ld_data_aligned_or_div[28]~q ),
	.prn(vcc));
defparam \av_ld_data_aligned_or_div[28] .is_wysiwyg = "true";
defparam \av_ld_data_aligned_or_div[28] .power_up = "low";

cyclonev_lcell_comb \E_stw_data[28]~26 (
	.dataa(!\E_src2_hazard_M~q ),
	.datab(!\M_ctrl_shift_rot~q ),
	.datac(!\av_ld_or_div_done~q ),
	.datad(!\M_shift_rot_result[28]~q ),
	.datae(!\av_ld_data_aligned_or_div[28]~q ),
	.dataf(!\M_alu_result[28]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_stw_data[28]~26_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_stw_data[28]~26 .extended_lut = "off";
defparam \E_stw_data[28]~26 .lut_mask = 64'h7DFFFFFFFFFFFFFF;
defparam \E_stw_data[28]~26 .shared_arith = "off";

cyclonev_lcell_comb \M_wr_data_unfiltered[28]~29 (
	.dataa(!\M_ctrl_shift_rot~q ),
	.datab(!\av_ld_or_div_done~q ),
	.datac(!\M_shift_rot_result[28]~q ),
	.datad(!\av_ld_data_aligned_or_div[28]~q ),
	.datae(!\M_alu_result[28]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_wr_data_unfiltered[28]~29_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_wr_data_unfiltered[28]~29 .extended_lut = "off";
defparam \M_wr_data_unfiltered[28]~29 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \M_wr_data_unfiltered[28]~29 .shared_arith = "off";

dffeas \W_wr_data[28] (
	.clk(clk_clk),
	.d(\M_wr_data_unfiltered[28]~29_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\W_wr_data[28]~q ),
	.prn(vcc));
defparam \W_wr_data[28] .is_wysiwyg = "true";
defparam \W_wr_data[28] .power_up = "low";

cyclonev_lcell_comb \D_src2_prelim[28]~24 (
	.dataa(!\M_wr_data_unfiltered[28]~29_combout ),
	.datab(!\D_src2_hazard_M~combout ),
	.datac(!\D_src2_hazard_W~combout ),
	.datad(!\W_wr_data[28]~q ),
	.datae(!\processor_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[28] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_prelim[28]~24_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_prelim[28]~24 .extended_lut = "off";
defparam \D_src2_prelim[28]~24 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \D_src2_prelim[28]~24 .shared_arith = "off";

dffeas \E_src2_prelim[28] (
	.clk(clk_clk),
	.d(\D_src2_prelim[28]~24_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_src2_prelim[28]~q ),
	.prn(vcc));
defparam \E_src2_prelim[28] .is_wysiwyg = "true";
defparam \E_src2_prelim[28] .power_up = "low";

cyclonev_lcell_comb \E_stw_data[28]~27 (
	.dataa(!\E_src2_hazard_M~q ),
	.datab(!\E_src2_prelim[28]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_stw_data[28]~27_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_stw_data[28]~27 .extended_lut = "off";
defparam \E_stw_data[28]~27 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \E_stw_data[28]~27 .shared_arith = "off";

cyclonev_lcell_comb \E_stw_data[28]~28 (
	.dataa(!\E_stw_data[28]~26_combout ),
	.datab(!\E_stw_data[28]~27_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_stw_data[28]~28_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_stw_data[28]~28 .extended_lut = "off";
defparam \E_stw_data[28]~28 .lut_mask = 64'h7777777777777777;
defparam \E_stw_data[28]~28 .shared_arith = "off";

dffeas \E_src2_imm[28] (
	.clk(clk_clk),
	.d(\D_iw[21]~q ),
	.asdata(\D_iw[18]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\D_ctrl_unsigned_lo_imm16~combout ),
	.sload(\Equal171~0_combout ),
	.ena(\W_stall~combout ),
	.q(\E_src2_imm[28]~q ),
	.prn(vcc));
defparam \E_src2_imm[28] .is_wysiwyg = "true";
defparam \E_src2_imm[28] .power_up = "low";

dffeas \d_readdata_d1[26] (
	.clk(clk_clk),
	.d(d_readdata[26]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d_readdata_d1[26]~q ),
	.prn(vcc));
defparam \d_readdata_d1[26] .is_wysiwyg = "true";
defparam \d_readdata_d1[26] .power_up = "low";

dffeas \av_ld_data_aligned_or_div[26] (
	.clk(clk_clk),
	.d(\av_fill_bit~0_combout ),
	.asdata(\d_readdata_d1[26]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\M_iw[4]~q ),
	.ena(vcc),
	.q(\av_ld_data_aligned_or_div[26]~q ),
	.prn(vcc));
defparam \av_ld_data_aligned_or_div[26] .is_wysiwyg = "true";
defparam \av_ld_data_aligned_or_div[26] .power_up = "low";

cyclonev_lcell_comb \E_stw_data[26]~38 (
	.dataa(!\E_src2_hazard_M~q ),
	.datab(!\M_ctrl_shift_rot~q ),
	.datac(!\av_ld_or_div_done~q ),
	.datad(!\M_shift_rot_result[26]~q ),
	.datae(!\av_ld_data_aligned_or_div[26]~q ),
	.dataf(!\M_alu_result[26]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_stw_data[26]~38_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_stw_data[26]~38 .extended_lut = "off";
defparam \E_stw_data[26]~38 .lut_mask = 64'h7DFFFFFFFFFFFFFF;
defparam \E_stw_data[26]~38 .shared_arith = "off";

cyclonev_lcell_comb \M_wr_data_unfiltered[26]~31 (
	.dataa(!\M_ctrl_shift_rot~q ),
	.datab(!\av_ld_or_div_done~q ),
	.datac(!\M_shift_rot_result[26]~q ),
	.datad(!\av_ld_data_aligned_or_div[26]~q ),
	.datae(!\M_alu_result[26]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_wr_data_unfiltered[26]~31_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_wr_data_unfiltered[26]~31 .extended_lut = "off";
defparam \M_wr_data_unfiltered[26]~31 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \M_wr_data_unfiltered[26]~31 .shared_arith = "off";

dffeas \W_wr_data[26] (
	.clk(clk_clk),
	.d(\M_wr_data_unfiltered[26]~31_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\W_wr_data[26]~q ),
	.prn(vcc));
defparam \W_wr_data[26] .is_wysiwyg = "true";
defparam \W_wr_data[26] .power_up = "low";

cyclonev_lcell_comb \D_src2_prelim[26]~29 (
	.dataa(!\M_wr_data_unfiltered[26]~31_combout ),
	.datab(!\D_src2_hazard_M~combout ),
	.datac(!\D_src2_hazard_W~combout ),
	.datad(!\W_wr_data[26]~q ),
	.datae(!\processor_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[26] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_prelim[26]~29_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_prelim[26]~29 .extended_lut = "off";
defparam \D_src2_prelim[26]~29 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \D_src2_prelim[26]~29 .shared_arith = "off";

dffeas \E_src2_prelim[26] (
	.clk(clk_clk),
	.d(\D_src2_prelim[26]~29_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_src2_prelim[26]~q ),
	.prn(vcc));
defparam \E_src2_prelim[26] .is_wysiwyg = "true";
defparam \E_src2_prelim[26] .power_up = "low";

cyclonev_lcell_comb \E_stw_data[26]~39 (
	.dataa(!\E_src2_hazard_M~q ),
	.datab(!\E_src2_prelim[26]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_stw_data[26]~39_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_stw_data[26]~39 .extended_lut = "off";
defparam \E_stw_data[26]~39 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \E_stw_data[26]~39 .shared_arith = "off";

cyclonev_lcell_comb \E_stw_data[26]~40 (
	.dataa(!\E_stw_data[26]~38_combout ),
	.datab(!\E_stw_data[26]~39_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_stw_data[26]~40_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_stw_data[26]~40 .extended_lut = "off";
defparam \E_stw_data[26]~40 .lut_mask = 64'h7777777777777777;
defparam \E_stw_data[26]~40 .shared_arith = "off";

dffeas \E_src2_imm[26] (
	.clk(clk_clk),
	.d(\D_iw[21]~q ),
	.asdata(\D_iw[16]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\D_ctrl_unsigned_lo_imm16~combout ),
	.sload(\Equal171~0_combout ),
	.ena(\W_stall~combout ),
	.q(\E_src2_imm[26]~q ),
	.prn(vcc));
defparam \E_src2_imm[26] .is_wysiwyg = "true";
defparam \E_src2_imm[26] .power_up = "low";

dffeas \d_readdata_d1[24] (
	.clk(clk_clk),
	.d(d_readdata[24]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d_readdata_d1[24]~q ),
	.prn(vcc));
defparam \d_readdata_d1[24] .is_wysiwyg = "true";
defparam \d_readdata_d1[24] .power_up = "low";

dffeas \av_ld_data_aligned_or_div[24] (
	.clk(clk_clk),
	.d(\av_fill_bit~0_combout ),
	.asdata(\d_readdata_d1[24]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\M_iw[4]~q ),
	.ena(vcc),
	.q(\av_ld_data_aligned_or_div[24]~q ),
	.prn(vcc));
defparam \av_ld_data_aligned_or_div[24] .is_wysiwyg = "true";
defparam \av_ld_data_aligned_or_div[24] .power_up = "low";

cyclonev_lcell_comb \E_stw_data[24]~18 (
	.dataa(!\E_src2_hazard_M~q ),
	.datab(!\M_ctrl_shift_rot~q ),
	.datac(!\av_ld_or_div_done~q ),
	.datad(!\M_shift_rot_result[24]~q ),
	.datae(!\av_ld_data_aligned_or_div[24]~q ),
	.dataf(!\M_alu_result[24]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_stw_data[24]~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_stw_data[24]~18 .extended_lut = "off";
defparam \E_stw_data[24]~18 .lut_mask = 64'h7DFFFFFFFFFFFFFF;
defparam \E_stw_data[24]~18 .shared_arith = "off";

cyclonev_lcell_comb \M_wr_data_unfiltered[24]~27 (
	.dataa(!\M_ctrl_shift_rot~q ),
	.datab(!\av_ld_or_div_done~q ),
	.datac(!\M_shift_rot_result[24]~q ),
	.datad(!\av_ld_data_aligned_or_div[24]~q ),
	.datae(!\M_alu_result[24]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_wr_data_unfiltered[24]~27_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_wr_data_unfiltered[24]~27 .extended_lut = "off";
defparam \M_wr_data_unfiltered[24]~27 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \M_wr_data_unfiltered[24]~27 .shared_arith = "off";

dffeas \W_wr_data[24] (
	.clk(clk_clk),
	.d(\M_wr_data_unfiltered[24]~27_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\W_wr_data[24]~q ),
	.prn(vcc));
defparam \W_wr_data[24] .is_wysiwyg = "true";
defparam \W_wr_data[24] .power_up = "low";

cyclonev_lcell_comb \D_src2_prelim[24]~20 (
	.dataa(!\M_wr_data_unfiltered[24]~27_combout ),
	.datab(!\D_src2_hazard_M~combout ),
	.datac(!\D_src2_hazard_W~combout ),
	.datad(!\W_wr_data[24]~q ),
	.datae(!\processor_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[24] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_prelim[24]~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_prelim[24]~20 .extended_lut = "off";
defparam \D_src2_prelim[24]~20 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \D_src2_prelim[24]~20 .shared_arith = "off";

dffeas \E_src2_prelim[24] (
	.clk(clk_clk),
	.d(\D_src2_prelim[24]~20_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_src2_prelim[24]~q ),
	.prn(vcc));
defparam \E_src2_prelim[24] .is_wysiwyg = "true";
defparam \E_src2_prelim[24] .power_up = "low";

cyclonev_lcell_comb \E_stw_data[24]~19 (
	.dataa(!\E_src2_hazard_M~q ),
	.datab(!\E_src2_prelim[24]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_stw_data[24]~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_stw_data[24]~19 .extended_lut = "off";
defparam \E_stw_data[24]~19 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \E_stw_data[24]~19 .shared_arith = "off";

cyclonev_lcell_comb \E_stw_data[24]~20 (
	.dataa(!\E_stw_data[24]~18_combout ),
	.datab(!\E_stw_data[24]~19_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_stw_data[24]~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_stw_data[24]~20 .extended_lut = "off";
defparam \E_stw_data[24]~20 .lut_mask = 64'h7777777777777777;
defparam \E_stw_data[24]~20 .shared_arith = "off";

dffeas \E_src2_imm[24] (
	.clk(clk_clk),
	.d(\D_iw[21]~q ),
	.asdata(\D_iw[14]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\D_ctrl_unsigned_lo_imm16~combout ),
	.sload(\Equal171~0_combout ),
	.ena(\W_stall~combout ),
	.q(\E_src2_imm[24]~q ),
	.prn(vcc));
defparam \E_src2_imm[24] .is_wysiwyg = "true";
defparam \E_src2_imm[24] .power_up = "low";

dffeas \d_readdata_d1[22] (
	.clk(clk_clk),
	.d(d_readdata[22]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d_readdata_d1[22]~q ),
	.prn(vcc));
defparam \d_readdata_d1[22] .is_wysiwyg = "true";
defparam \d_readdata_d1[22] .power_up = "low";

dffeas \av_ld_data_aligned_or_div[22] (
	.clk(clk_clk),
	.d(\av_fill_bit~0_combout ),
	.asdata(\d_readdata_d1[22]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\M_iw[4]~q ),
	.ena(vcc),
	.q(\av_ld_data_aligned_or_div[22]~q ),
	.prn(vcc));
defparam \av_ld_data_aligned_or_div[22] .is_wysiwyg = "true";
defparam \av_ld_data_aligned_or_div[22] .power_up = "low";

cyclonev_lcell_comb \E_stw_data[22]~29 (
	.dataa(!\E_src2_hazard_M~q ),
	.datab(!\M_ctrl_shift_rot~q ),
	.datac(!\av_ld_or_div_done~q ),
	.datad(!\M_shift_rot_result[22]~q ),
	.datae(!\av_ld_data_aligned_or_div[22]~q ),
	.dataf(!\M_alu_result[22]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_stw_data[22]~29_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_stw_data[22]~29 .extended_lut = "off";
defparam \E_stw_data[22]~29 .lut_mask = 64'h7DFFFFFFFFFFFFFF;
defparam \E_stw_data[22]~29 .shared_arith = "off";

cyclonev_lcell_comb \M_wr_data_unfiltered[22]~30 (
	.dataa(!\M_ctrl_shift_rot~q ),
	.datab(!\av_ld_or_div_done~q ),
	.datac(!\M_shift_rot_result[22]~q ),
	.datad(!\av_ld_data_aligned_or_div[22]~q ),
	.datae(!\M_alu_result[22]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_wr_data_unfiltered[22]~30_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_wr_data_unfiltered[22]~30 .extended_lut = "off";
defparam \M_wr_data_unfiltered[22]~30 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \M_wr_data_unfiltered[22]~30 .shared_arith = "off";

dffeas \W_wr_data[22] (
	.clk(clk_clk),
	.d(\M_wr_data_unfiltered[22]~30_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\W_wr_data[22]~q ),
	.prn(vcc));
defparam \W_wr_data[22] .is_wysiwyg = "true";
defparam \W_wr_data[22] .power_up = "low";

cyclonev_lcell_comb \D_src2_prelim[22]~25 (
	.dataa(!\M_wr_data_unfiltered[22]~30_combout ),
	.datab(!\D_src2_hazard_M~combout ),
	.datac(!\D_src2_hazard_W~combout ),
	.datad(!\W_wr_data[22]~q ),
	.datae(!\processor_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[22] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_prelim[22]~25_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_prelim[22]~25 .extended_lut = "off";
defparam \D_src2_prelim[22]~25 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \D_src2_prelim[22]~25 .shared_arith = "off";

dffeas \E_src2_prelim[22] (
	.clk(clk_clk),
	.d(\D_src2_prelim[22]~25_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_src2_prelim[22]~q ),
	.prn(vcc));
defparam \E_src2_prelim[22] .is_wysiwyg = "true";
defparam \E_src2_prelim[22] .power_up = "low";

cyclonev_lcell_comb \E_stw_data[22]~30 (
	.dataa(!\E_src2_hazard_M~q ),
	.datab(!\E_src2_prelim[22]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_stw_data[22]~30_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_stw_data[22]~30 .extended_lut = "off";
defparam \E_stw_data[22]~30 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \E_stw_data[22]~30 .shared_arith = "off";

cyclonev_lcell_comb \E_stw_data[22]~31 (
	.dataa(!\E_stw_data[22]~29_combout ),
	.datab(!\E_stw_data[22]~30_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_stw_data[22]~31_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_stw_data[22]~31 .extended_lut = "off";
defparam \E_stw_data[22]~31 .lut_mask = 64'h7777777777777777;
defparam \E_stw_data[22]~31 .shared_arith = "off";

dffeas \E_src2_imm[22] (
	.clk(clk_clk),
	.d(\D_iw[21]~q ),
	.asdata(\D_iw[12]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\D_ctrl_unsigned_lo_imm16~combout ),
	.sload(\Equal171~0_combout ),
	.ena(\W_stall~combout ),
	.q(\E_src2_imm[22]~q ),
	.prn(vcc));
defparam \E_src2_imm[22] .is_wysiwyg = "true";
defparam \E_src2_imm[22] .power_up = "low";

dffeas \d_readdata_d1[20] (
	.clk(clk_clk),
	.d(d_readdata[20]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d_readdata_d1[20]~q ),
	.prn(vcc));
defparam \d_readdata_d1[20] .is_wysiwyg = "true";
defparam \d_readdata_d1[20] .power_up = "low";

dffeas \av_ld_data_aligned_or_div[20] (
	.clk(clk_clk),
	.d(\av_fill_bit~0_combout ),
	.asdata(\d_readdata_d1[20]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\M_iw[4]~q ),
	.ena(vcc),
	.q(\av_ld_data_aligned_or_div[20]~q ),
	.prn(vcc));
defparam \av_ld_data_aligned_or_div[20] .is_wysiwyg = "true";
defparam \av_ld_data_aligned_or_div[20] .power_up = "low";

cyclonev_lcell_comb \E_stw_data[20]~23 (
	.dataa(!\E_src2_hazard_M~q ),
	.datab(!\M_ctrl_shift_rot~q ),
	.datac(!\av_ld_or_div_done~q ),
	.datad(!\M_shift_rot_result[20]~q ),
	.datae(!\av_ld_data_aligned_or_div[20]~q ),
	.dataf(!\M_alu_result[20]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_stw_data[20]~23_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_stw_data[20]~23 .extended_lut = "off";
defparam \E_stw_data[20]~23 .lut_mask = 64'h7DFFFFFFFFFFFFFF;
defparam \E_stw_data[20]~23 .shared_arith = "off";

cyclonev_lcell_comb \M_wr_data_unfiltered[20]~28 (
	.dataa(!\M_ctrl_shift_rot~q ),
	.datab(!\av_ld_or_div_done~q ),
	.datac(!\M_shift_rot_result[20]~q ),
	.datad(!\av_ld_data_aligned_or_div[20]~q ),
	.datae(!\M_alu_result[20]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_wr_data_unfiltered[20]~28_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_wr_data_unfiltered[20]~28 .extended_lut = "off";
defparam \M_wr_data_unfiltered[20]~28 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \M_wr_data_unfiltered[20]~28 .shared_arith = "off";

dffeas \W_wr_data[20] (
	.clk(clk_clk),
	.d(\M_wr_data_unfiltered[20]~28_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\W_wr_data[20]~q ),
	.prn(vcc));
defparam \W_wr_data[20] .is_wysiwyg = "true";
defparam \W_wr_data[20] .power_up = "low";

cyclonev_lcell_comb \D_src2_prelim[20]~23 (
	.dataa(!\M_wr_data_unfiltered[20]~28_combout ),
	.datab(!\D_src2_hazard_M~combout ),
	.datac(!\D_src2_hazard_W~combout ),
	.datad(!\W_wr_data[20]~q ),
	.datae(!\processor_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[20] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_prelim[20]~23_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_prelim[20]~23 .extended_lut = "off";
defparam \D_src2_prelim[20]~23 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \D_src2_prelim[20]~23 .shared_arith = "off";

dffeas \E_src2_prelim[20] (
	.clk(clk_clk),
	.d(\D_src2_prelim[20]~23_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_src2_prelim[20]~q ),
	.prn(vcc));
defparam \E_src2_prelim[20] .is_wysiwyg = "true";
defparam \E_src2_prelim[20] .power_up = "low";

cyclonev_lcell_comb \E_stw_data[20]~24 (
	.dataa(!\E_src2_hazard_M~q ),
	.datab(!\E_src2_prelim[20]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_stw_data[20]~24_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_stw_data[20]~24 .extended_lut = "off";
defparam \E_stw_data[20]~24 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \E_stw_data[20]~24 .shared_arith = "off";

cyclonev_lcell_comb \E_stw_data[20]~25 (
	.dataa(!\E_stw_data[20]~23_combout ),
	.datab(!\E_stw_data[20]~24_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_stw_data[20]~25_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_stw_data[20]~25 .extended_lut = "off";
defparam \E_stw_data[20]~25 .lut_mask = 64'h7777777777777777;
defparam \E_stw_data[20]~25 .shared_arith = "off";

cyclonev_lcell_comb \F_iw[10]~24 (
	.dataa(!\intr_req~0_combout ),
	.datab(!\processor_cpu_ic_data|the_altsyncram|auto_generated|q_b[10] ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[10]~24_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[10]~24 .extended_lut = "off";
defparam \F_iw[10]~24 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \F_iw[10]~24 .shared_arith = "off";

dffeas \D_iw[10] (
	.clk(clk_clk),
	.d(\F_iw[10]~24_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\F_iw~1_combout ),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\D_iw[10]~q ),
	.prn(vcc));
defparam \D_iw[10] .is_wysiwyg = "true";
defparam \D_iw[10] .power_up = "low";

dffeas \E_src2_imm[20] (
	.clk(clk_clk),
	.d(\D_iw[21]~q ),
	.asdata(\D_iw[10]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\D_ctrl_unsigned_lo_imm16~combout ),
	.sload(\Equal171~0_combout ),
	.ena(\W_stall~combout ),
	.q(\E_src2_imm[20]~q ),
	.prn(vcc));
defparam \E_src2_imm[20] .is_wysiwyg = "true";
defparam \E_src2_imm[20] .power_up = "low";

dffeas \d_readdata_d1[18] (
	.clk(clk_clk),
	.d(d_readdata[18]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d_readdata_d1[18]~q ),
	.prn(vcc));
defparam \d_readdata_d1[18] .is_wysiwyg = "true";
defparam \d_readdata_d1[18] .power_up = "low";

dffeas \av_ld_data_aligned_or_div[18] (
	.clk(clk_clk),
	.d(\av_fill_bit~0_combout ),
	.asdata(\d_readdata_d1[18]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\M_iw[4]~q ),
	.ena(vcc),
	.q(\av_ld_data_aligned_or_div[18]~q ),
	.prn(vcc));
defparam \av_ld_data_aligned_or_div[18] .is_wysiwyg = "true";
defparam \av_ld_data_aligned_or_div[18] .power_up = "low";

cyclonev_lcell_comb \E_stw_data[18]~32 (
	.dataa(!\E_src2_hazard_M~q ),
	.datab(!\M_ctrl_shift_rot~q ),
	.datac(!\av_ld_or_div_done~q ),
	.datad(!\M_shift_rot_result[18]~q ),
	.datae(!\av_ld_data_aligned_or_div[18]~q ),
	.dataf(!\M_alu_result[18]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_stw_data[18]~32_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_stw_data[18]~32 .extended_lut = "off";
defparam \E_stw_data[18]~32 .lut_mask = 64'h7DFFFFFFFFFFFFFF;
defparam \E_stw_data[18]~32 .shared_arith = "off";

cyclonev_lcell_comb \M_wr_data_unfiltered[18]~23 (
	.dataa(!\M_ctrl_shift_rot~q ),
	.datab(!\av_ld_or_div_done~q ),
	.datac(!\M_shift_rot_result[18]~q ),
	.datad(!\av_ld_data_aligned_or_div[18]~q ),
	.datae(!\M_alu_result[18]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_wr_data_unfiltered[18]~23_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_wr_data_unfiltered[18]~23 .extended_lut = "off";
defparam \M_wr_data_unfiltered[18]~23 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \M_wr_data_unfiltered[18]~23 .shared_arith = "off";

dffeas \W_wr_data[18] (
	.clk(clk_clk),
	.d(\M_wr_data_unfiltered[18]~23_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\W_wr_data[18]~q ),
	.prn(vcc));
defparam \W_wr_data[18] .is_wysiwyg = "true";
defparam \W_wr_data[18] .power_up = "low";

cyclonev_lcell_comb \D_src2_prelim[18]~26 (
	.dataa(!\M_wr_data_unfiltered[18]~23_combout ),
	.datab(!\D_src2_hazard_M~combout ),
	.datac(!\D_src2_hazard_W~combout ),
	.datad(!\W_wr_data[18]~q ),
	.datae(!\processor_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[18] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_prelim[18]~26_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_prelim[18]~26 .extended_lut = "off";
defparam \D_src2_prelim[18]~26 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \D_src2_prelim[18]~26 .shared_arith = "off";

dffeas \E_src2_prelim[18] (
	.clk(clk_clk),
	.d(\D_src2_prelim[18]~26_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_src2_prelim[18]~q ),
	.prn(vcc));
defparam \E_src2_prelim[18] .is_wysiwyg = "true";
defparam \E_src2_prelim[18] .power_up = "low";

cyclonev_lcell_comb \E_stw_data[18]~33 (
	.dataa(!\E_src2_hazard_M~q ),
	.datab(!\E_src2_prelim[18]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_stw_data[18]~33_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_stw_data[18]~33 .extended_lut = "off";
defparam \E_stw_data[18]~33 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \E_stw_data[18]~33 .shared_arith = "off";

cyclonev_lcell_comb \E_stw_data[18]~34 (
	.dataa(!\E_stw_data[18]~32_combout ),
	.datab(!\E_stw_data[18]~33_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_stw_data[18]~34_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_stw_data[18]~34 .extended_lut = "off";
defparam \E_stw_data[18]~34 .lut_mask = 64'h7777777777777777;
defparam \E_stw_data[18]~34 .shared_arith = "off";

cyclonev_lcell_comb \F_iw[8]~26 (
	.dataa(!\intr_req~0_combout ),
	.datab(!\processor_cpu_ic_data|the_altsyncram|auto_generated|q_b[8] ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[8]~26_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[8]~26 .extended_lut = "off";
defparam \F_iw[8]~26 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \F_iw[8]~26 .shared_arith = "off";

dffeas \D_iw[8] (
	.clk(clk_clk),
	.d(\F_iw[8]~26_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\F_iw~1_combout ),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\D_iw[8]~q ),
	.prn(vcc));
defparam \D_iw[8] .is_wysiwyg = "true";
defparam \D_iw[8] .power_up = "low";

dffeas \E_src2_imm[18] (
	.clk(clk_clk),
	.d(\D_iw[21]~q ),
	.asdata(\D_iw[8]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\D_ctrl_unsigned_lo_imm16~combout ),
	.sload(\Equal171~0_combout ),
	.ena(\W_stall~combout ),
	.q(\E_src2_imm[18]~q ),
	.prn(vcc));
defparam \E_src2_imm[18] .is_wysiwyg = "true";
defparam \E_src2_imm[18] .power_up = "low";

dffeas \d_readdata_d1[16] (
	.clk(clk_clk),
	.d(d_readdata[16]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d_readdata_d1[16]~q ),
	.prn(vcc));
defparam \d_readdata_d1[16] .is_wysiwyg = "true";
defparam \d_readdata_d1[16] .power_up = "low";

dffeas \av_ld_data_aligned_or_div[16] (
	.clk(clk_clk),
	.d(\av_fill_bit~0_combout ),
	.asdata(\d_readdata_d1[16]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\M_iw[4]~q ),
	.ena(vcc),
	.q(\av_ld_data_aligned_or_div[16]~q ),
	.prn(vcc));
defparam \av_ld_data_aligned_or_div[16] .is_wysiwyg = "true";
defparam \av_ld_data_aligned_or_div[16] .power_up = "low";

cyclonev_lcell_comb \E_src1[16]~7 (
	.dataa(!M_alu_result_16),
	.datab(!\M_ctrl_shift_rot~q ),
	.datac(!\av_ld_or_div_done~q ),
	.datad(!\E_src1_hazard_M~q ),
	.datae(!\M_shift_rot_result[16]~q ),
	.dataf(!\av_ld_data_aligned_or_div[16]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_src1[16]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_src1[16]~7 .extended_lut = "off";
defparam \E_src1[16]~7 .lut_mask = 64'h7DFFFFFFFFFFFFFF;
defparam \E_src1[16]~7 .shared_arith = "off";

cyclonev_lcell_comb \M_wr_data_unfiltered[16]~13 (
	.dataa(!M_alu_result_16),
	.datab(!\M_ctrl_shift_rot~q ),
	.datac(!\av_ld_or_div_done~q ),
	.datad(!\M_shift_rot_result[16]~q ),
	.datae(!\av_ld_data_aligned_or_div[16]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_wr_data_unfiltered[16]~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_wr_data_unfiltered[16]~13 .extended_lut = "off";
defparam \M_wr_data_unfiltered[16]~13 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \M_wr_data_unfiltered[16]~13 .shared_arith = "off";

cyclonev_lcell_comb \D_src1_hazard_M~0 (
	.dataa(!\M_wr_dst_reg~q ),
	.datab(!\M_dst_regnum[0]~q ),
	.datac(!\M_dst_regnum[1]~q ),
	.datad(!\D_iw[27]~q ),
	.datae(!\D_iw[28]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_hazard_M~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src1_hazard_M~0 .extended_lut = "off";
defparam \D_src1_hazard_M~0 .lut_mask = 64'hBEEBEBBEBEEBEBBE;
defparam \D_src1_hazard_M~0 .shared_arith = "off";

cyclonev_lcell_comb \D_src1_hazard_M~1 (
	.dataa(!\M_dst_regnum[2]~q ),
	.datab(!\M_dst_regnum[3]~q ),
	.datac(!\D_iw[29]~q ),
	.datad(!\D_iw[30]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_hazard_M~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src1_hazard_M~1 .extended_lut = "off";
defparam \D_src1_hazard_M~1 .lut_mask = 64'h6996699669966996;
defparam \D_src1_hazard_M~1 .shared_arith = "off";

cyclonev_lcell_comb D_src1_hazard_M(
	.dataa(!\M_dst_regnum[4]~q ),
	.datab(!\D_ctrl_a_not_src~0_combout ),
	.datac(!\D_iw[31]~q ),
	.datad(!\D_src1_hazard_M~0_combout ),
	.datae(!\D_src1_hazard_M~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_hazard_M~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam D_src1_hazard_M.extended_lut = "off";
defparam D_src1_hazard_M.lut_mask = 64'hDEFFFFFFDEFFFFFF;
defparam D_src1_hazard_M.shared_arith = "off";

cyclonev_lcell_comb \D_src1_hazard_W~0 (
	.dataa(!\W_wr_dst_reg~q ),
	.datab(!\W_dst_regnum[0]~q ),
	.datac(!\W_dst_regnum[1]~q ),
	.datad(!\D_iw[27]~q ),
	.datae(!\D_iw[28]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_hazard_W~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src1_hazard_W~0 .extended_lut = "off";
defparam \D_src1_hazard_W~0 .lut_mask = 64'h7DD7D77D7DD7D77D;
defparam \D_src1_hazard_W~0 .shared_arith = "off";

cyclonev_lcell_comb \D_src1_hazard_W~1 (
	.dataa(!\W_dst_regnum[2]~q ),
	.datab(!\W_dst_regnum[3]~q ),
	.datac(!\D_iw[29]~q ),
	.datad(!\D_iw[30]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_hazard_W~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src1_hazard_W~1 .extended_lut = "off";
defparam \D_src1_hazard_W~1 .lut_mask = 64'h6996699669966996;
defparam \D_src1_hazard_W~1 .shared_arith = "off";

cyclonev_lcell_comb D_src1_hazard_W(
	.dataa(!\W_dst_regnum[4]~q ),
	.datab(!\D_ctrl_a_not_src~0_combout ),
	.datac(!\D_iw[31]~q ),
	.datad(!\D_src1_hazard_W~0_combout ),
	.datae(!\D_src1_hazard_W~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_hazard_W~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam D_src1_hazard_W.extended_lut = "off";
defparam D_src1_hazard_W.lut_mask = 64'hDEFFFFFFDEFFFFFF;
defparam D_src1_hazard_W.shared_arith = "off";

dffeas \W_wr_data[16] (
	.clk(clk_clk),
	.d(\M_wr_data_unfiltered[16]~13_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\W_wr_data[16]~q ),
	.prn(vcc));
defparam \W_wr_data[16] .is_wysiwyg = "true";
defparam \W_wr_data[16] .power_up = "low";

cyclonev_lcell_comb \D_src1_prelim[16]~3 (
	.dataa(!\M_wr_data_unfiltered[16]~13_combout ),
	.datab(!\D_src1_hazard_M~combout ),
	.datac(!\D_src1_hazard_W~combout ),
	.datad(!\W_wr_data[16]~q ),
	.datae(!\processor_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[16] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_prelim[16]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src1_prelim[16]~3 .extended_lut = "off";
defparam \D_src1_prelim[16]~3 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \D_src1_prelim[16]~3 .shared_arith = "off";

dffeas \E_src1_prelim[16] (
	.clk(clk_clk),
	.d(\D_src1_prelim[16]~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_src1_prelim[16]~q ),
	.prn(vcc));
defparam \E_src1_prelim[16] .is_wysiwyg = "true";
defparam \E_src1_prelim[16] .power_up = "low";

cyclonev_lcell_comb \E_src1[16]~8 (
	.dataa(!\E_src1_hazard_M~q ),
	.datab(!\E_src1_prelim[16]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_src1[16]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_src1[16]~8 .extended_lut = "off";
defparam \E_src1[16]~8 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \E_src1[16]~8 .shared_arith = "off";

cyclonev_lcell_comb \E_src1[16]~9 (
	.dataa(!\E_src1[16]~7_combout ),
	.datab(!\E_src1[16]~8_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_src1[16]~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_src1[16]~9 .extended_lut = "off";
defparam \E_src1[16]~9 .lut_mask = 64'h7777777777777777;
defparam \E_src1[16]~9 .shared_arith = "off";

cyclonev_lcell_comb \Equal2~0 (
	.dataa(!\M_iw[4]~q ),
	.datab(!\M_iw[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal2~0 .extended_lut = "off";
defparam \Equal2~0 .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \Equal2~0 .shared_arith = "off";

cyclonev_lcell_comb \av_ld_byte1_data[7]~0 (
	.dataa(!\M_ld_align_sh16~combout ),
	.datab(!\Equal2~0_combout ),
	.datac(!\d_readdata_d1[15]~q ),
	.datad(!\d_readdata_d1[31]~q ),
	.datae(!\av_fill_bit~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_ld_byte1_data[7]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_ld_byte1_data[7]~0 .extended_lut = "off";
defparam \av_ld_byte1_data[7]~0 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \av_ld_byte1_data[7]~0 .shared_arith = "off";

dffeas \av_ld_data_aligned_or_div[15] (
	.clk(clk_clk),
	.d(\av_ld_byte1_data[7]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\av_ld_data_aligned_or_div[15]~q ),
	.prn(vcc));
defparam \av_ld_data_aligned_or_div[15] .is_wysiwyg = "true";
defparam \av_ld_data_aligned_or_div[15] .power_up = "low";

cyclonev_lcell_comb \M_wr_data_unfiltered[15]~1 (
	.dataa(!M_alu_result_15),
	.datab(!\M_ctrl_shift_rot~q ),
	.datac(!\av_ld_or_div_done~q ),
	.datad(!\M_shift_rot_result[15]~q ),
	.datae(!\av_ld_data_aligned_or_div[15]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_wr_data_unfiltered[15]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_wr_data_unfiltered[15]~1 .extended_lut = "off";
defparam \M_wr_data_unfiltered[15]~1 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \M_wr_data_unfiltered[15]~1 .shared_arith = "off";

dffeas \W_wr_data[15] (
	.clk(clk_clk),
	.d(\M_wr_data_unfiltered[15]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\W_wr_data[15]~q ),
	.prn(vcc));
defparam \W_wr_data[15] .is_wysiwyg = "true";
defparam \W_wr_data[15] .power_up = "low";

cyclonev_lcell_comb \D_src1_prelim[15]~4 (
	.dataa(!\M_wr_data_unfiltered[15]~1_combout ),
	.datab(!\D_src1_hazard_M~combout ),
	.datac(!\D_src1_hazard_W~combout ),
	.datad(!\W_wr_data[15]~q ),
	.datae(!\processor_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[15] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_prelim[15]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src1_prelim[15]~4 .extended_lut = "off";
defparam \D_src1_prelim[15]~4 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \D_src1_prelim[15]~4 .shared_arith = "off";

dffeas \E_src1_prelim[15] (
	.clk(clk_clk),
	.d(\D_src1_prelim[15]~4_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_src1_prelim[15]~q ),
	.prn(vcc));
defparam \E_src1_prelim[15] .is_wysiwyg = "true";
defparam \E_src1_prelim[15] .power_up = "low";

cyclonev_lcell_comb \E_src1[15]~10 (
	.dataa(!\E_src1_hazard_M~q ),
	.datab(!\M_wr_data_unfiltered[15]~1_combout ),
	.datac(!\E_src1_prelim[15]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_src1[15]~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_src1[15]~10 .extended_lut = "off";
defparam \E_src1[15]~10 .lut_mask = 64'h2727272727272727;
defparam \E_src1[15]~10 .shared_arith = "off";

dffeas \d_readdata_d1[14] (
	.clk(clk_clk),
	.d(d_readdata[14]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d_readdata_d1[14]~q ),
	.prn(vcc));
defparam \d_readdata_d1[14] .is_wysiwyg = "true";
defparam \d_readdata_d1[14] .power_up = "low";

cyclonev_lcell_comb \av_ld_byte1_data[6]~1 (
	.dataa(!\M_ld_align_sh16~combout ),
	.datab(!\Equal2~0_combout ),
	.datac(!\d_readdata_d1[14]~q ),
	.datad(!\d_readdata_d1[30]~q ),
	.datae(!\av_fill_bit~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_ld_byte1_data[6]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_ld_byte1_data[6]~1 .extended_lut = "off";
defparam \av_ld_byte1_data[6]~1 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \av_ld_byte1_data[6]~1 .shared_arith = "off";

dffeas \av_ld_data_aligned_or_div[14] (
	.clk(clk_clk),
	.d(\av_ld_byte1_data[6]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\av_ld_data_aligned_or_div[14]~q ),
	.prn(vcc));
defparam \av_ld_data_aligned_or_div[14] .is_wysiwyg = "true";
defparam \av_ld_data_aligned_or_div[14] .power_up = "low";

cyclonev_lcell_comb \M_wr_data_unfiltered[14]~2 (
	.dataa(!M_alu_result_14),
	.datab(!\M_ctrl_shift_rot~q ),
	.datac(!\av_ld_or_div_done~q ),
	.datad(!\M_shift_rot_result[14]~q ),
	.datae(!\av_ld_data_aligned_or_div[14]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_wr_data_unfiltered[14]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_wr_data_unfiltered[14]~2 .extended_lut = "off";
defparam \M_wr_data_unfiltered[14]~2 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \M_wr_data_unfiltered[14]~2 .shared_arith = "off";

dffeas \W_wr_data[14] (
	.clk(clk_clk),
	.d(\M_wr_data_unfiltered[14]~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\W_wr_data[14]~q ),
	.prn(vcc));
defparam \W_wr_data[14] .is_wysiwyg = "true";
defparam \W_wr_data[14] .power_up = "low";

cyclonev_lcell_comb \D_src1_prelim[14]~5 (
	.dataa(!\M_wr_data_unfiltered[14]~2_combout ),
	.datab(!\D_src1_hazard_M~combout ),
	.datac(!\D_src1_hazard_W~combout ),
	.datad(!\W_wr_data[14]~q ),
	.datae(!\processor_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[14] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_prelim[14]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src1_prelim[14]~5 .extended_lut = "off";
defparam \D_src1_prelim[14]~5 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \D_src1_prelim[14]~5 .shared_arith = "off";

dffeas \E_src1_prelim[14] (
	.clk(clk_clk),
	.d(\D_src1_prelim[14]~5_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_src1_prelim[14]~q ),
	.prn(vcc));
defparam \E_src1_prelim[14] .is_wysiwyg = "true";
defparam \E_src1_prelim[14] .power_up = "low";

cyclonev_lcell_comb \E_src1[14]~11 (
	.dataa(!\E_src1_hazard_M~q ),
	.datab(!\M_wr_data_unfiltered[14]~2_combout ),
	.datac(!\E_src1_prelim[14]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_src1[14]~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_src1[14]~11 .extended_lut = "off";
defparam \E_src1[14]~11 .lut_mask = 64'h2727272727272727;
defparam \E_src1[14]~11 .shared_arith = "off";

dffeas \d_readdata_d1[12] (
	.clk(clk_clk),
	.d(d_readdata[12]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d_readdata_d1[12]~q ),
	.prn(vcc));
defparam \d_readdata_d1[12] .is_wysiwyg = "true";
defparam \d_readdata_d1[12] .power_up = "low";

cyclonev_lcell_comb \av_ld_byte1_data[4]~3 (
	.dataa(!\M_ld_align_sh16~combout ),
	.datab(!\Equal2~0_combout ),
	.datac(!\d_readdata_d1[12]~q ),
	.datad(!\d_readdata_d1[28]~q ),
	.datae(!\av_fill_bit~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_ld_byte1_data[4]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_ld_byte1_data[4]~3 .extended_lut = "off";
defparam \av_ld_byte1_data[4]~3 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \av_ld_byte1_data[4]~3 .shared_arith = "off";

dffeas \av_ld_data_aligned_or_div[12] (
	.clk(clk_clk),
	.d(\av_ld_byte1_data[4]~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\av_ld_data_aligned_or_div[12]~q ),
	.prn(vcc));
defparam \av_ld_data_aligned_or_div[12] .is_wysiwyg = "true";
defparam \av_ld_data_aligned_or_div[12] .power_up = "low";

cyclonev_lcell_comb \M_wr_data_unfiltered[12]~4 (
	.dataa(!M_alu_result_12),
	.datab(!\M_ctrl_shift_rot~q ),
	.datac(!\av_ld_or_div_done~q ),
	.datad(!\M_shift_rot_result[12]~q ),
	.datae(!\av_ld_data_aligned_or_div[12]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_wr_data_unfiltered[12]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_wr_data_unfiltered[12]~4 .extended_lut = "off";
defparam \M_wr_data_unfiltered[12]~4 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \M_wr_data_unfiltered[12]~4 .shared_arith = "off";

dffeas \W_wr_data[12] (
	.clk(clk_clk),
	.d(\M_wr_data_unfiltered[12]~4_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\W_wr_data[12]~q ),
	.prn(vcc));
defparam \W_wr_data[12] .is_wysiwyg = "true";
defparam \W_wr_data[12] .power_up = "low";

cyclonev_lcell_comb \D_src1_prelim[12]~7 (
	.dataa(!\M_wr_data_unfiltered[12]~4_combout ),
	.datab(!\D_src1_hazard_M~combout ),
	.datac(!\D_src1_hazard_W~combout ),
	.datad(!\W_wr_data[12]~q ),
	.datae(!\processor_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[12] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_prelim[12]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src1_prelim[12]~7 .extended_lut = "off";
defparam \D_src1_prelim[12]~7 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \D_src1_prelim[12]~7 .shared_arith = "off";

dffeas \E_src1_prelim[12] (
	.clk(clk_clk),
	.d(\D_src1_prelim[12]~7_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_src1_prelim[12]~q ),
	.prn(vcc));
defparam \E_src1_prelim[12] .is_wysiwyg = "true";
defparam \E_src1_prelim[12] .power_up = "low";

cyclonev_lcell_comb \E_src1[12]~13 (
	.dataa(!\E_src1_hazard_M~q ),
	.datab(!\M_wr_data_unfiltered[12]~4_combout ),
	.datac(!\E_src1_prelim[12]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_src1[12]~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_src1[12]~13 .extended_lut = "off";
defparam \E_src1[12]~13 .lut_mask = 64'h2727272727272727;
defparam \E_src1[12]~13 .shared_arith = "off";

cyclonev_lcell_comb \av_ld_byte1_data[3]~4 (
	.dataa(!\M_ld_align_sh16~combout ),
	.datab(!\Equal2~0_combout ),
	.datac(!\d_readdata_d1[11]~q ),
	.datad(!\d_readdata_d1[27]~q ),
	.datae(!\av_fill_bit~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_ld_byte1_data[3]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_ld_byte1_data[3]~4 .extended_lut = "off";
defparam \av_ld_byte1_data[3]~4 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \av_ld_byte1_data[3]~4 .shared_arith = "off";

dffeas \av_ld_data_aligned_or_div[11] (
	.clk(clk_clk),
	.d(\av_ld_byte1_data[3]~4_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\av_ld_data_aligned_or_div[11]~q ),
	.prn(vcc));
defparam \av_ld_data_aligned_or_div[11] .is_wysiwyg = "true";
defparam \av_ld_data_aligned_or_div[11] .power_up = "low";

cyclonev_lcell_comb \M_wr_data_unfiltered[11]~5 (
	.dataa(!M_alu_result_11),
	.datab(!\M_ctrl_shift_rot~q ),
	.datac(!\av_ld_or_div_done~q ),
	.datad(!\M_shift_rot_result[11]~q ),
	.datae(!\av_ld_data_aligned_or_div[11]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_wr_data_unfiltered[11]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_wr_data_unfiltered[11]~5 .extended_lut = "off";
defparam \M_wr_data_unfiltered[11]~5 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \M_wr_data_unfiltered[11]~5 .shared_arith = "off";

dffeas \W_wr_data[11] (
	.clk(clk_clk),
	.d(\M_wr_data_unfiltered[11]~5_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\W_wr_data[11]~q ),
	.prn(vcc));
defparam \W_wr_data[11] .is_wysiwyg = "true";
defparam \W_wr_data[11] .power_up = "low";

cyclonev_lcell_comb \D_src1_prelim[11]~8 (
	.dataa(!\M_wr_data_unfiltered[11]~5_combout ),
	.datab(!\D_src1_hazard_M~combout ),
	.datac(!\D_src1_hazard_W~combout ),
	.datad(!\W_wr_data[11]~q ),
	.datae(!\processor_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[11] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_prelim[11]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src1_prelim[11]~8 .extended_lut = "off";
defparam \D_src1_prelim[11]~8 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \D_src1_prelim[11]~8 .shared_arith = "off";

dffeas \E_src1_prelim[11] (
	.clk(clk_clk),
	.d(\D_src1_prelim[11]~8_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_src1_prelim[11]~q ),
	.prn(vcc));
defparam \E_src1_prelim[11] .is_wysiwyg = "true";
defparam \E_src1_prelim[11] .power_up = "low";

cyclonev_lcell_comb \E_src1[11]~14 (
	.dataa(!\E_src1_hazard_M~q ),
	.datab(!\M_wr_data_unfiltered[11]~5_combout ),
	.datac(!\E_src1_prelim[11]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_src1[11]~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_src1[11]~14 .extended_lut = "off";
defparam \E_src1[11]~14 .lut_mask = 64'h2727272727272727;
defparam \E_src1[11]~14 .shared_arith = "off";

dffeas \d_readdata_d1[10] (
	.clk(clk_clk),
	.d(d_readdata[10]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d_readdata_d1[10]~q ),
	.prn(vcc));
defparam \d_readdata_d1[10] .is_wysiwyg = "true";
defparam \d_readdata_d1[10] .power_up = "low";

cyclonev_lcell_comb \av_ld_byte1_data[2]~5 (
	.dataa(!\M_ld_align_sh16~combout ),
	.datab(!\Equal2~0_combout ),
	.datac(!\d_readdata_d1[10]~q ),
	.datad(!\d_readdata_d1[26]~q ),
	.datae(!\av_fill_bit~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_ld_byte1_data[2]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_ld_byte1_data[2]~5 .extended_lut = "off";
defparam \av_ld_byte1_data[2]~5 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \av_ld_byte1_data[2]~5 .shared_arith = "off";

dffeas \av_ld_data_aligned_or_div[10] (
	.clk(clk_clk),
	.d(\av_ld_byte1_data[2]~5_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\av_ld_data_aligned_or_div[10]~q ),
	.prn(vcc));
defparam \av_ld_data_aligned_or_div[10] .is_wysiwyg = "true";
defparam \av_ld_data_aligned_or_div[10] .power_up = "low";

cyclonev_lcell_comb \E_src1[10]~15 (
	.dataa(!M_alu_result_10),
	.datab(!\M_ctrl_shift_rot~q ),
	.datac(!\av_ld_or_div_done~q ),
	.datad(!\E_src1_hazard_M~q ),
	.datae(!\M_shift_rot_result[10]~q ),
	.dataf(!\av_ld_data_aligned_or_div[10]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_src1[10]~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_src1[10]~15 .extended_lut = "off";
defparam \E_src1[10]~15 .lut_mask = 64'h7DFFFFFFFFFFFFFF;
defparam \E_src1[10]~15 .shared_arith = "off";

cyclonev_lcell_comb \M_wr_data_unfiltered[10]~14 (
	.dataa(!M_alu_result_10),
	.datab(!\M_ctrl_shift_rot~q ),
	.datac(!\av_ld_or_div_done~q ),
	.datad(!\M_shift_rot_result[10]~q ),
	.datae(!\av_ld_data_aligned_or_div[10]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_wr_data_unfiltered[10]~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_wr_data_unfiltered[10]~14 .extended_lut = "off";
defparam \M_wr_data_unfiltered[10]~14 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \M_wr_data_unfiltered[10]~14 .shared_arith = "off";

dffeas \W_wr_data[10] (
	.clk(clk_clk),
	.d(\M_wr_data_unfiltered[10]~14_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\W_wr_data[10]~q ),
	.prn(vcc));
defparam \W_wr_data[10] .is_wysiwyg = "true";
defparam \W_wr_data[10] .power_up = "low";

cyclonev_lcell_comb \D_src1_prelim[10]~9 (
	.dataa(!\M_wr_data_unfiltered[10]~14_combout ),
	.datab(!\D_src1_hazard_M~combout ),
	.datac(!\D_src1_hazard_W~combout ),
	.datad(!\W_wr_data[10]~q ),
	.datae(!\processor_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[10] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_prelim[10]~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src1_prelim[10]~9 .extended_lut = "off";
defparam \D_src1_prelim[10]~9 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \D_src1_prelim[10]~9 .shared_arith = "off";

dffeas \E_src1_prelim[10] (
	.clk(clk_clk),
	.d(\D_src1_prelim[10]~9_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_src1_prelim[10]~q ),
	.prn(vcc));
defparam \E_src1_prelim[10] .is_wysiwyg = "true";
defparam \E_src1_prelim[10] .power_up = "low";

cyclonev_lcell_comb \E_src1[10]~16 (
	.dataa(!\E_src1_hazard_M~q ),
	.datab(!\E_src1_prelim[10]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_src1[10]~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_src1[10]~16 .extended_lut = "off";
defparam \E_src1[10]~16 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \E_src1[10]~16 .shared_arith = "off";

cyclonev_lcell_comb \E_src1[10]~17 (
	.dataa(!\E_src1[10]~15_combout ),
	.datab(!\E_src1[10]~16_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_src1[10]~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_src1[10]~17 .extended_lut = "off";
defparam \E_src1[10]~17 .lut_mask = 64'h7777777777777777;
defparam \E_src1[10]~17 .shared_arith = "off";

cyclonev_lcell_comb \av_ld_byte1_data[1]~6 (
	.dataa(!\M_ld_align_sh16~combout ),
	.datab(!\Equal2~0_combout ),
	.datac(!\av_fill_bit~0_combout ),
	.datad(!\d_readdata_d1[25]~q ),
	.datae(!\d_readdata_d1[9]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_ld_byte1_data[1]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_ld_byte1_data[1]~6 .extended_lut = "off";
defparam \av_ld_byte1_data[1]~6 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \av_ld_byte1_data[1]~6 .shared_arith = "off";

dffeas \av_ld_data_aligned_or_div[9] (
	.clk(clk_clk),
	.d(\av_ld_byte1_data[1]~6_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\av_ld_data_aligned_or_div[9]~q ),
	.prn(vcc));
defparam \av_ld_data_aligned_or_div[9] .is_wysiwyg = "true";
defparam \av_ld_data_aligned_or_div[9] .power_up = "low";

cyclonev_lcell_comb \M_wr_data_unfiltered[9]~6 (
	.dataa(!M_alu_result_9),
	.datab(!\M_ctrl_shift_rot~q ),
	.datac(!\av_ld_or_div_done~q ),
	.datad(!\M_shift_rot_result[9]~q ),
	.datae(!\av_ld_data_aligned_or_div[9]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_wr_data_unfiltered[9]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_wr_data_unfiltered[9]~6 .extended_lut = "off";
defparam \M_wr_data_unfiltered[9]~6 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \M_wr_data_unfiltered[9]~6 .shared_arith = "off";

dffeas \W_wr_data[9] (
	.clk(clk_clk),
	.d(\M_wr_data_unfiltered[9]~6_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\W_wr_data[9]~q ),
	.prn(vcc));
defparam \W_wr_data[9] .is_wysiwyg = "true";
defparam \W_wr_data[9] .power_up = "low";

cyclonev_lcell_comb \D_src1_prelim[9]~10 (
	.dataa(!\M_wr_data_unfiltered[9]~6_combout ),
	.datab(!\D_src1_hazard_M~combout ),
	.datac(!\D_src1_hazard_W~combout ),
	.datad(!\W_wr_data[9]~q ),
	.datae(!\processor_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[9] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_prelim[9]~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src1_prelim[9]~10 .extended_lut = "off";
defparam \D_src1_prelim[9]~10 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \D_src1_prelim[9]~10 .shared_arith = "off";

dffeas \E_src1_prelim[9] (
	.clk(clk_clk),
	.d(\D_src1_prelim[9]~10_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_src1_prelim[9]~q ),
	.prn(vcc));
defparam \E_src1_prelim[9] .is_wysiwyg = "true";
defparam \E_src1_prelim[9] .power_up = "low";

cyclonev_lcell_comb \E_src1[9]~18 (
	.dataa(!\E_src1_hazard_M~q ),
	.datab(!\M_wr_data_unfiltered[9]~6_combout ),
	.datac(!\E_src1_prelim[9]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_src1[9]~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_src1[9]~18 .extended_lut = "off";
defparam \E_src1[9]~18 .lut_mask = 64'h2727272727272727;
defparam \E_src1[9]~18 .shared_arith = "off";

dffeas \d_readdata_d1[8] (
	.clk(clk_clk),
	.d(d_readdata[8]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d_readdata_d1[8]~q ),
	.prn(vcc));
defparam \d_readdata_d1[8] .is_wysiwyg = "true";
defparam \d_readdata_d1[8] .power_up = "low";

cyclonev_lcell_comb \av_ld_byte1_data[0]~7 (
	.dataa(!\d_readdata_d1[8]~q ),
	.datab(!\d_readdata_d1[24]~q ),
	.datac(!\M_ld_align_sh16~combout ),
	.datad(!\Equal2~0_combout ),
	.datae(!\av_fill_bit~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_ld_byte1_data[0]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_ld_byte1_data[0]~7 .extended_lut = "off";
defparam \av_ld_byte1_data[0]~7 .lut_mask = 64'h7FF7FFFF7FF7FFFF;
defparam \av_ld_byte1_data[0]~7 .shared_arith = "off";

dffeas \av_ld_data_aligned_or_div[8] (
	.clk(clk_clk),
	.d(\av_ld_byte1_data[0]~7_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\av_ld_data_aligned_or_div[8]~q ),
	.prn(vcc));
defparam \av_ld_data_aligned_or_div[8] .is_wysiwyg = "true";
defparam \av_ld_data_aligned_or_div[8] .power_up = "low";

cyclonev_lcell_comb \E_src1[8]~19 (
	.dataa(!M_alu_result_8),
	.datab(!\M_ctrl_shift_rot~q ),
	.datac(!\av_ld_or_div_done~q ),
	.datad(!\E_src1_hazard_M~q ),
	.datae(!\M_shift_rot_result[8]~q ),
	.dataf(!\av_ld_data_aligned_or_div[8]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_src1[8]~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_src1[8]~19 .extended_lut = "off";
defparam \E_src1[8]~19 .lut_mask = 64'h7DFFFFFFFFFFFFFF;
defparam \E_src1[8]~19 .shared_arith = "off";

cyclonev_lcell_comb \M_wr_data_unfiltered[8]~15 (
	.dataa(!M_alu_result_8),
	.datab(!\M_ctrl_shift_rot~q ),
	.datac(!\av_ld_or_div_done~q ),
	.datad(!\M_shift_rot_result[8]~q ),
	.datae(!\av_ld_data_aligned_or_div[8]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_wr_data_unfiltered[8]~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_wr_data_unfiltered[8]~15 .extended_lut = "off";
defparam \M_wr_data_unfiltered[8]~15 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \M_wr_data_unfiltered[8]~15 .shared_arith = "off";

dffeas \W_wr_data[8] (
	.clk(clk_clk),
	.d(\M_wr_data_unfiltered[8]~15_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\W_wr_data[8]~q ),
	.prn(vcc));
defparam \W_wr_data[8] .is_wysiwyg = "true";
defparam \W_wr_data[8] .power_up = "low";

cyclonev_lcell_comb \D_src1_prelim[8]~11 (
	.dataa(!\M_wr_data_unfiltered[8]~15_combout ),
	.datab(!\D_src1_hazard_M~combout ),
	.datac(!\D_src1_hazard_W~combout ),
	.datad(!\W_wr_data[8]~q ),
	.datae(!\processor_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[8] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_prelim[8]~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src1_prelim[8]~11 .extended_lut = "off";
defparam \D_src1_prelim[8]~11 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \D_src1_prelim[8]~11 .shared_arith = "off";

dffeas \E_src1_prelim[8] (
	.clk(clk_clk),
	.d(\D_src1_prelim[8]~11_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_src1_prelim[8]~q ),
	.prn(vcc));
defparam \E_src1_prelim[8] .is_wysiwyg = "true";
defparam \E_src1_prelim[8] .power_up = "low";

cyclonev_lcell_comb \E_src1[8]~20 (
	.dataa(!\E_src1_hazard_M~q ),
	.datab(!\E_src1_prelim[8]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_src1[8]~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_src1[8]~20 .extended_lut = "off";
defparam \E_src1[8]~20 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \E_src1[8]~20 .shared_arith = "off";

cyclonev_lcell_comb \E_src1[8]~21 (
	.dataa(!\E_src1[8]~19_combout ),
	.datab(!\E_src1[8]~20_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_src1[8]~21_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_src1[8]~21 .extended_lut = "off";
defparam \E_src1[8]~21 .lut_mask = 64'h7777777777777777;
defparam \E_src1[8]~21 .shared_arith = "off";

dffeas \d_readdata_d1[5] (
	.clk(clk_clk),
	.d(d_readdata[5]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d_readdata_d1[5]~q ),
	.prn(vcc));
defparam \d_readdata_d1[5] .is_wysiwyg = "true";
defparam \d_readdata_d1[5] .power_up = "low";

dffeas \d_readdata_d1[21] (
	.clk(clk_clk),
	.d(d_readdata[21]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d_readdata_d1[21]~q ),
	.prn(vcc));
defparam \d_readdata_d1[21] .is_wysiwyg = "true";
defparam \d_readdata_d1[21] .power_up = "low";

dffeas \d_readdata_d1[13] (
	.clk(clk_clk),
	.d(d_readdata[13]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d_readdata_d1[13]~q ),
	.prn(vcc));
defparam \d_readdata_d1[13] .is_wysiwyg = "true";
defparam \d_readdata_d1[13] .power_up = "low";

dffeas \d_readdata_d1[29] (
	.clk(clk_clk),
	.d(d_readdata[29]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d_readdata_d1[29]~q ),
	.prn(vcc));
defparam \d_readdata_d1[29] .is_wysiwyg = "true";
defparam \d_readdata_d1[29] .power_up = "low";

cyclonev_lcell_comb \av_ld_byte0_data[5]~1 (
	.dataa(!\d_readdata_d1[5]~q ),
	.datab(!\d_readdata_d1[21]~q ),
	.datac(!\d_readdata_d1[13]~q ),
	.datad(!\d_readdata_d1[29]~q ),
	.datae(!\M_ld_align_sh16~combout ),
	.dataf(!\M_ld_align_sh8~combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_ld_byte0_data[5]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_ld_byte0_data[5]~1 .extended_lut = "off";
defparam \av_ld_byte0_data[5]~1 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \av_ld_byte0_data[5]~1 .shared_arith = "off";

dffeas \av_ld_data_aligned_or_div[5] (
	.clk(clk_clk),
	.d(\av_ld_byte0_data[5]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\av_ld_data_aligned_or_div[5]~q ),
	.prn(vcc));
defparam \av_ld_data_aligned_or_div[5] .is_wysiwyg = "true";
defparam \av_ld_data_aligned_or_div[5] .power_up = "low";

cyclonev_lcell_comb \M_wr_data_unfiltered[5]~0 (
	.dataa(!M_alu_result_5),
	.datab(!\M_ctrl_shift_rot~q ),
	.datac(!\av_ld_or_div_done~q ),
	.datad(!\M_shift_rot_result[5]~q ),
	.datae(!\av_ld_data_aligned_or_div[5]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_wr_data_unfiltered[5]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_wr_data_unfiltered[5]~0 .extended_lut = "off";
defparam \M_wr_data_unfiltered[5]~0 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \M_wr_data_unfiltered[5]~0 .shared_arith = "off";

dffeas \W_wr_data[5] (
	.clk(clk_clk),
	.d(\M_wr_data_unfiltered[5]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\W_wr_data[5]~q ),
	.prn(vcc));
defparam \W_wr_data[5] .is_wysiwyg = "true";
defparam \W_wr_data[5] .power_up = "low";

cyclonev_lcell_comb \D_src1_prelim[5]~0 (
	.dataa(!\M_wr_data_unfiltered[5]~0_combout ),
	.datab(!\D_src1_hazard_M~combout ),
	.datac(!\D_src1_hazard_W~combout ),
	.datad(!\W_wr_data[5]~q ),
	.datae(!\processor_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[5] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_prelim[5]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src1_prelim[5]~0 .extended_lut = "off";
defparam \D_src1_prelim[5]~0 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \D_src1_prelim[5]~0 .shared_arith = "off";

dffeas \E_src1_prelim[5] (
	.clk(clk_clk),
	.d(\D_src1_prelim[5]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_src1_prelim[5]~q ),
	.prn(vcc));
defparam \E_src1_prelim[5] .is_wysiwyg = "true";
defparam \E_src1_prelim[5] .power_up = "low";

cyclonev_lcell_comb \E_src1[5]~0 (
	.dataa(!\E_src1_hazard_M~q ),
	.datab(!\M_wr_data_unfiltered[5]~0_combout ),
	.datac(!\E_src1_prelim[5]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_src1[5]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_src1[5]~0 .extended_lut = "off";
defparam \E_src1[5]~0 .lut_mask = 64'h2727272727272727;
defparam \E_src1[5]~0 .shared_arith = "off";

dffeas \d_readdata_d1[4] (
	.clk(clk_clk),
	.d(d_readdata[4]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d_readdata_d1[4]~q ),
	.prn(vcc));
defparam \d_readdata_d1[4] .is_wysiwyg = "true";
defparam \d_readdata_d1[4] .power_up = "low";

cyclonev_lcell_comb \av_ld_byte0_data[4]~2 (
	.dataa(!\d_readdata_d1[4]~q ),
	.datab(!\d_readdata_d1[20]~q ),
	.datac(!\d_readdata_d1[12]~q ),
	.datad(!\d_readdata_d1[28]~q ),
	.datae(!\M_ld_align_sh16~combout ),
	.dataf(!\M_ld_align_sh8~combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_ld_byte0_data[4]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_ld_byte0_data[4]~2 .extended_lut = "off";
defparam \av_ld_byte0_data[4]~2 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \av_ld_byte0_data[4]~2 .shared_arith = "off";

dffeas \av_ld_data_aligned_or_div[4] (
	.clk(clk_clk),
	.d(\av_ld_byte0_data[4]~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\av_ld_data_aligned_or_div[4]~q ),
	.prn(vcc));
defparam \av_ld_data_aligned_or_div[4] .is_wysiwyg = "true";
defparam \av_ld_data_aligned_or_div[4] .power_up = "low";

cyclonev_lcell_comb \E_src1[4]~1 (
	.dataa(!M_alu_result_4),
	.datab(!\M_ctrl_shift_rot~q ),
	.datac(!\av_ld_or_div_done~q ),
	.datad(!\E_src1_hazard_M~q ),
	.datae(!\M_shift_rot_result[4]~q ),
	.dataf(!\av_ld_data_aligned_or_div[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_src1[4]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_src1[4]~1 .extended_lut = "off";
defparam \E_src1[4]~1 .lut_mask = 64'h7DFFFFFFFFFFFFFF;
defparam \E_src1[4]~1 .shared_arith = "off";

cyclonev_lcell_comb \M_wr_data_unfiltered[4]~11 (
	.dataa(!M_alu_result_4),
	.datab(!\M_ctrl_shift_rot~q ),
	.datac(!\av_ld_or_div_done~q ),
	.datad(!\M_shift_rot_result[4]~q ),
	.datae(!\av_ld_data_aligned_or_div[4]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_wr_data_unfiltered[4]~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_wr_data_unfiltered[4]~11 .extended_lut = "off";
defparam \M_wr_data_unfiltered[4]~11 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \M_wr_data_unfiltered[4]~11 .shared_arith = "off";

dffeas \W_wr_data[4] (
	.clk(clk_clk),
	.d(\M_wr_data_unfiltered[4]~11_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\W_wr_data[4]~q ),
	.prn(vcc));
defparam \W_wr_data[4] .is_wysiwyg = "true";
defparam \W_wr_data[4] .power_up = "low";

cyclonev_lcell_comb \D_src1_prelim[4]~1 (
	.dataa(!\M_wr_data_unfiltered[4]~11_combout ),
	.datab(!\D_src1_hazard_M~combout ),
	.datac(!\D_src1_hazard_W~combout ),
	.datad(!\W_wr_data[4]~q ),
	.datae(!\processor_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[4] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_prelim[4]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src1_prelim[4]~1 .extended_lut = "off";
defparam \D_src1_prelim[4]~1 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \D_src1_prelim[4]~1 .shared_arith = "off";

dffeas \E_src1_prelim[4] (
	.clk(clk_clk),
	.d(\D_src1_prelim[4]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_src1_prelim[4]~q ),
	.prn(vcc));
defparam \E_src1_prelim[4] .is_wysiwyg = "true";
defparam \E_src1_prelim[4] .power_up = "low";

cyclonev_lcell_comb \E_src1[4]~2 (
	.dataa(!\E_src1_hazard_M~q ),
	.datab(!\E_src1_prelim[4]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_src1[4]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_src1[4]~2 .extended_lut = "off";
defparam \E_src1[4]~2 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \E_src1[4]~2 .shared_arith = "off";

cyclonev_lcell_comb \E_src1[4]~3 (
	.dataa(!\E_src1[4]~1_combout ),
	.datab(!\E_src1[4]~2_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_src1[4]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_src1[4]~3 .extended_lut = "off";
defparam \E_src1[4]~3 .lut_mask = 64'h7777777777777777;
defparam \E_src1[4]~3 .shared_arith = "off";

cyclonev_lcell_comb \M_shift_rot_result_nxt[4]~2 (
	.dataa(!\M_shift_rot_stall~q ),
	.datab(!\M_shift_rot_result[3]~q ),
	.datac(!\M_shift_rot_result[5]~q ),
	.datad(!\E_src1[4]~3_combout ),
	.datae(!\M_ctrl_shift_rot_right~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_shift_rot_result_nxt[4]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_shift_rot_result_nxt[4]~2 .extended_lut = "off";
defparam \M_shift_rot_result_nxt[4]~2 .lut_mask = 64'h7FFFBFFF7FFFBFFF;
defparam \M_shift_rot_result_nxt[4]~2 .shared_arith = "off";

dffeas \M_shift_rot_result[4] (
	.clk(clk_clk),
	.d(\M_shift_rot_result_nxt[4]~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\M_shift_rot_result[4]~q ),
	.prn(vcc));
defparam \M_shift_rot_result[4] .is_wysiwyg = "true";
defparam \M_shift_rot_result[4] .power_up = "low";

cyclonev_lcell_comb \M_shift_rot_result_nxt[5]~1 (
	.dataa(!\M_shift_rot_stall~q ),
	.datab(!\E_src1[5]~0_combout ),
	.datac(!\M_shift_rot_result[4]~q ),
	.datad(!\M_shift_rot_result[6]~q ),
	.datae(!\M_ctrl_shift_rot_right~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_shift_rot_result_nxt[5]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_shift_rot_result_nxt[5]~1 .extended_lut = "off";
defparam \M_shift_rot_result_nxt[5]~1 .lut_mask = 64'h7FFFBFFF7FFFBFFF;
defparam \M_shift_rot_result_nxt[5]~1 .shared_arith = "off";

dffeas \M_shift_rot_result[5] (
	.clk(clk_clk),
	.d(\M_shift_rot_result_nxt[5]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\M_shift_rot_result[5]~q ),
	.prn(vcc));
defparam \M_shift_rot_result[5] .is_wysiwyg = "true";
defparam \M_shift_rot_result[5] .power_up = "low";

dffeas \d_readdata_d1[6] (
	.clk(clk_clk),
	.d(d_readdata[6]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d_readdata_d1[6]~q ),
	.prn(vcc));
defparam \d_readdata_d1[6] .is_wysiwyg = "true";
defparam \d_readdata_d1[6] .power_up = "low";

cyclonev_lcell_comb \av_ld_byte0_data[6]~3 (
	.dataa(!\d_readdata_d1[6]~q ),
	.datab(!\d_readdata_d1[22]~q ),
	.datac(!\d_readdata_d1[14]~q ),
	.datad(!\d_readdata_d1[30]~q ),
	.datae(!\M_ld_align_sh16~combout ),
	.dataf(!\M_ld_align_sh8~combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_ld_byte0_data[6]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_ld_byte0_data[6]~3 .extended_lut = "off";
defparam \av_ld_byte0_data[6]~3 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \av_ld_byte0_data[6]~3 .shared_arith = "off";

dffeas \av_ld_data_aligned_or_div[6] (
	.clk(clk_clk),
	.d(\av_ld_byte0_data[6]~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\av_ld_data_aligned_or_div[6]~q ),
	.prn(vcc));
defparam \av_ld_data_aligned_or_div[6] .is_wysiwyg = "true";
defparam \av_ld_data_aligned_or_div[6] .power_up = "low";

cyclonev_lcell_comb \E_src1[6]~4 (
	.dataa(!M_alu_result_6),
	.datab(!\M_ctrl_shift_rot~q ),
	.datac(!\av_ld_or_div_done~q ),
	.datad(!\E_src1_hazard_M~q ),
	.datae(!\M_shift_rot_result[6]~q ),
	.dataf(!\av_ld_data_aligned_or_div[6]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_src1[6]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_src1[6]~4 .extended_lut = "off";
defparam \E_src1[6]~4 .lut_mask = 64'h7DFFFFFFFFFFFFFF;
defparam \E_src1[6]~4 .shared_arith = "off";

cyclonev_lcell_comb \M_wr_data_unfiltered[6]~12 (
	.dataa(!M_alu_result_6),
	.datab(!\M_ctrl_shift_rot~q ),
	.datac(!\av_ld_or_div_done~q ),
	.datad(!\M_shift_rot_result[6]~q ),
	.datae(!\av_ld_data_aligned_or_div[6]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_wr_data_unfiltered[6]~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_wr_data_unfiltered[6]~12 .extended_lut = "off";
defparam \M_wr_data_unfiltered[6]~12 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \M_wr_data_unfiltered[6]~12 .shared_arith = "off";

dffeas \W_wr_data[6] (
	.clk(clk_clk),
	.d(\M_wr_data_unfiltered[6]~12_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\W_wr_data[6]~q ),
	.prn(vcc));
defparam \W_wr_data[6] .is_wysiwyg = "true";
defparam \W_wr_data[6] .power_up = "low";

cyclonev_lcell_comb \D_src1_prelim[6]~2 (
	.dataa(!\M_wr_data_unfiltered[6]~12_combout ),
	.datab(!\D_src1_hazard_M~combout ),
	.datac(!\D_src1_hazard_W~combout ),
	.datad(!\W_wr_data[6]~q ),
	.datae(!\processor_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[6] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_prelim[6]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src1_prelim[6]~2 .extended_lut = "off";
defparam \D_src1_prelim[6]~2 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \D_src1_prelim[6]~2 .shared_arith = "off";

dffeas \E_src1_prelim[6] (
	.clk(clk_clk),
	.d(\D_src1_prelim[6]~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_src1_prelim[6]~q ),
	.prn(vcc));
defparam \E_src1_prelim[6] .is_wysiwyg = "true";
defparam \E_src1_prelim[6] .power_up = "low";

cyclonev_lcell_comb \E_src1[6]~5 (
	.dataa(!\E_src1_hazard_M~q ),
	.datab(!\E_src1_prelim[6]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_src1[6]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_src1[6]~5 .extended_lut = "off";
defparam \E_src1[6]~5 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \E_src1[6]~5 .shared_arith = "off";

cyclonev_lcell_comb \E_src1[6]~6 (
	.dataa(!\E_src1[6]~4_combout ),
	.datab(!\E_src1[6]~5_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_src1[6]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_src1[6]~6 .extended_lut = "off";
defparam \E_src1[6]~6 .lut_mask = 64'h7777777777777777;
defparam \E_src1[6]~6 .shared_arith = "off";

cyclonev_lcell_comb \M_shift_rot_result_nxt[6]~3 (
	.dataa(!\M_shift_rot_stall~q ),
	.datab(!\M_shift_rot_result[5]~q ),
	.datac(!\E_src1[6]~6_combout ),
	.datad(!\M_shift_rot_result[7]~q ),
	.datae(!\M_ctrl_shift_rot_right~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_shift_rot_result_nxt[6]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_shift_rot_result_nxt[6]~3 .extended_lut = "off";
defparam \M_shift_rot_result_nxt[6]~3 .lut_mask = 64'h7FFFBFFF7FFFBFFF;
defparam \M_shift_rot_result_nxt[6]~3 .shared_arith = "off";

dffeas \M_shift_rot_result[6] (
	.clk(clk_clk),
	.d(\M_shift_rot_result_nxt[6]~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\M_shift_rot_result[6]~q ),
	.prn(vcc));
defparam \M_shift_rot_result[6] .is_wysiwyg = "true";
defparam \M_shift_rot_result[6] .power_up = "low";

cyclonev_lcell_comb \av_ld_byte0_data[7]~4 (
	.dataa(!\d_readdata_d1[7]~q ),
	.datab(!\d_readdata_d1[23]~q ),
	.datac(!\d_readdata_d1[15]~q ),
	.datad(!\d_readdata_d1[31]~q ),
	.datae(!\M_ld_align_sh16~combout ),
	.dataf(!\M_ld_align_sh8~combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_ld_byte0_data[7]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_ld_byte0_data[7]~4 .extended_lut = "off";
defparam \av_ld_byte0_data[7]~4 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \av_ld_byte0_data[7]~4 .shared_arith = "off";

dffeas \av_ld_data_aligned_or_div[7] (
	.clk(clk_clk),
	.d(\av_ld_byte0_data[7]~4_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\av_ld_data_aligned_or_div[7]~q ),
	.prn(vcc));
defparam \av_ld_data_aligned_or_div[7] .is_wysiwyg = "true";
defparam \av_ld_data_aligned_or_div[7] .power_up = "low";

cyclonev_lcell_comb \M_wr_data_unfiltered[7]~7 (
	.dataa(!M_alu_result_7),
	.datab(!\M_ctrl_shift_rot~q ),
	.datac(!\av_ld_or_div_done~q ),
	.datad(!\M_shift_rot_result[7]~q ),
	.datae(!\av_ld_data_aligned_or_div[7]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_wr_data_unfiltered[7]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_wr_data_unfiltered[7]~7 .extended_lut = "off";
defparam \M_wr_data_unfiltered[7]~7 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \M_wr_data_unfiltered[7]~7 .shared_arith = "off";

dffeas \W_wr_data[7] (
	.clk(clk_clk),
	.d(\M_wr_data_unfiltered[7]~7_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\W_wr_data[7]~q ),
	.prn(vcc));
defparam \W_wr_data[7] .is_wysiwyg = "true";
defparam \W_wr_data[7] .power_up = "low";

cyclonev_lcell_comb \D_src1_prelim[7]~12 (
	.dataa(!\M_wr_data_unfiltered[7]~7_combout ),
	.datab(!\D_src1_hazard_M~combout ),
	.datac(!\D_src1_hazard_W~combout ),
	.datad(!\W_wr_data[7]~q ),
	.datae(!\processor_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[7] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_prelim[7]~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src1_prelim[7]~12 .extended_lut = "off";
defparam \D_src1_prelim[7]~12 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \D_src1_prelim[7]~12 .shared_arith = "off";

dffeas \E_src1_prelim[7] (
	.clk(clk_clk),
	.d(\D_src1_prelim[7]~12_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_src1_prelim[7]~q ),
	.prn(vcc));
defparam \E_src1_prelim[7] .is_wysiwyg = "true";
defparam \E_src1_prelim[7] .power_up = "low";

cyclonev_lcell_comb \E_src1[7]~22 (
	.dataa(!\E_src1_hazard_M~q ),
	.datab(!\M_wr_data_unfiltered[7]~7_combout ),
	.datac(!\E_src1_prelim[7]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_src1[7]~22_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_src1[7]~22 .extended_lut = "off";
defparam \E_src1[7]~22 .lut_mask = 64'h2727272727272727;
defparam \E_src1[7]~22 .shared_arith = "off";

cyclonev_lcell_comb \M_shift_rot_result_nxt[7]~13 (
	.dataa(!\M_shift_rot_stall~q ),
	.datab(!\M_shift_rot_result[6]~q ),
	.datac(!\M_shift_rot_result[8]~q ),
	.datad(!\E_src1[7]~22_combout ),
	.datae(!\M_ctrl_shift_rot_right~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_shift_rot_result_nxt[7]~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_shift_rot_result_nxt[7]~13 .extended_lut = "off";
defparam \M_shift_rot_result_nxt[7]~13 .lut_mask = 64'h7FFFBFFF7FFFBFFF;
defparam \M_shift_rot_result_nxt[7]~13 .shared_arith = "off";

dffeas \M_shift_rot_result[7] (
	.clk(clk_clk),
	.d(\M_shift_rot_result_nxt[7]~13_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\M_shift_rot_result[7]~q ),
	.prn(vcc));
defparam \M_shift_rot_result[7] .is_wysiwyg = "true";
defparam \M_shift_rot_result[7] .power_up = "low";

cyclonev_lcell_comb \M_shift_rot_result_nxt[8]~12 (
	.dataa(!\M_shift_rot_stall~q ),
	.datab(!\M_shift_rot_result[9]~q ),
	.datac(!\E_src1[8]~21_combout ),
	.datad(!\M_shift_rot_result[7]~q ),
	.datae(!\M_ctrl_shift_rot_right~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_shift_rot_result_nxt[8]~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_shift_rot_result_nxt[8]~12 .extended_lut = "off";
defparam \M_shift_rot_result_nxt[8]~12 .lut_mask = 64'h7FFFBFFF7FFFBFFF;
defparam \M_shift_rot_result_nxt[8]~12 .shared_arith = "off";

dffeas \M_shift_rot_result[8] (
	.clk(clk_clk),
	.d(\M_shift_rot_result_nxt[8]~12_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\M_shift_rot_result[8]~q ),
	.prn(vcc));
defparam \M_shift_rot_result[8] .is_wysiwyg = "true";
defparam \M_shift_rot_result[8] .power_up = "low";

cyclonev_lcell_comb \M_shift_rot_result_nxt[9]~11 (
	.dataa(!\M_shift_rot_stall~q ),
	.datab(!\M_shift_rot_result[10]~q ),
	.datac(!\E_src1[9]~18_combout ),
	.datad(!\M_shift_rot_result[8]~q ),
	.datae(!\M_ctrl_shift_rot_right~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_shift_rot_result_nxt[9]~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_shift_rot_result_nxt[9]~11 .extended_lut = "off";
defparam \M_shift_rot_result_nxt[9]~11 .lut_mask = 64'h7FFFBFFF7FFFBFFF;
defparam \M_shift_rot_result_nxt[9]~11 .shared_arith = "off";

dffeas \M_shift_rot_result[9] (
	.clk(clk_clk),
	.d(\M_shift_rot_result_nxt[9]~11_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\M_shift_rot_result[9]~q ),
	.prn(vcc));
defparam \M_shift_rot_result[9] .is_wysiwyg = "true";
defparam \M_shift_rot_result[9] .power_up = "low";

cyclonev_lcell_comb \M_shift_rot_result_nxt[10]~10 (
	.dataa(!\M_shift_rot_stall~q ),
	.datab(!\M_shift_rot_result[11]~q ),
	.datac(!\E_src1[10]~17_combout ),
	.datad(!\M_shift_rot_result[9]~q ),
	.datae(!\M_ctrl_shift_rot_right~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_shift_rot_result_nxt[10]~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_shift_rot_result_nxt[10]~10 .extended_lut = "off";
defparam \M_shift_rot_result_nxt[10]~10 .lut_mask = 64'h7FFFBFFF7FFFBFFF;
defparam \M_shift_rot_result_nxt[10]~10 .shared_arith = "off";

dffeas \M_shift_rot_result[10] (
	.clk(clk_clk),
	.d(\M_shift_rot_result_nxt[10]~10_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\M_shift_rot_result[10]~q ),
	.prn(vcc));
defparam \M_shift_rot_result[10] .is_wysiwyg = "true";
defparam \M_shift_rot_result[10] .power_up = "low";

cyclonev_lcell_comb \M_shift_rot_result_nxt[11]~9 (
	.dataa(!\M_shift_rot_stall~q ),
	.datab(!\M_shift_rot_result[12]~q ),
	.datac(!\E_src1[11]~14_combout ),
	.datad(!\M_shift_rot_result[10]~q ),
	.datae(!\M_ctrl_shift_rot_right~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_shift_rot_result_nxt[11]~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_shift_rot_result_nxt[11]~9 .extended_lut = "off";
defparam \M_shift_rot_result_nxt[11]~9 .lut_mask = 64'h7FFFBFFF7FFFBFFF;
defparam \M_shift_rot_result_nxt[11]~9 .shared_arith = "off";

dffeas \M_shift_rot_result[11] (
	.clk(clk_clk),
	.d(\M_shift_rot_result_nxt[11]~9_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\M_shift_rot_result[11]~q ),
	.prn(vcc));
defparam \M_shift_rot_result[11] .is_wysiwyg = "true";
defparam \M_shift_rot_result[11] .power_up = "low";

cyclonev_lcell_comb \M_shift_rot_result_nxt[12]~8 (
	.dataa(!\M_shift_rot_stall~q ),
	.datab(!\E_src1[12]~13_combout ),
	.datac(!\M_shift_rot_result[11]~q ),
	.datad(!\M_shift_rot_result[13]~q ),
	.datae(!\M_ctrl_shift_rot_right~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_shift_rot_result_nxt[12]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_shift_rot_result_nxt[12]~8 .extended_lut = "off";
defparam \M_shift_rot_result_nxt[12]~8 .lut_mask = 64'h7FFFBFFF7FFFBFFF;
defparam \M_shift_rot_result_nxt[12]~8 .shared_arith = "off";

dffeas \M_shift_rot_result[12] (
	.clk(clk_clk),
	.d(\M_shift_rot_result_nxt[12]~8_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\M_shift_rot_result[12]~q ),
	.prn(vcc));
defparam \M_shift_rot_result[12] .is_wysiwyg = "true";
defparam \M_shift_rot_result[12] .power_up = "low";

cyclonev_lcell_comb \av_ld_byte1_data[5]~2 (
	.dataa(!\M_ld_align_sh16~combout ),
	.datab(!\Equal2~0_combout ),
	.datac(!\d_readdata_d1[13]~q ),
	.datad(!\d_readdata_d1[29]~q ),
	.datae(!\av_fill_bit~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_ld_byte1_data[5]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_ld_byte1_data[5]~2 .extended_lut = "off";
defparam \av_ld_byte1_data[5]~2 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \av_ld_byte1_data[5]~2 .shared_arith = "off";

dffeas \av_ld_data_aligned_or_div[13] (
	.clk(clk_clk),
	.d(\av_ld_byte1_data[5]~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\av_ld_data_aligned_or_div[13]~q ),
	.prn(vcc));
defparam \av_ld_data_aligned_or_div[13] .is_wysiwyg = "true";
defparam \av_ld_data_aligned_or_div[13] .power_up = "low";

cyclonev_lcell_comb \M_wr_data_unfiltered[13]~3 (
	.dataa(!M_alu_result_13),
	.datab(!\M_ctrl_shift_rot~q ),
	.datac(!\av_ld_or_div_done~q ),
	.datad(!\M_shift_rot_result[13]~q ),
	.datae(!\av_ld_data_aligned_or_div[13]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_wr_data_unfiltered[13]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_wr_data_unfiltered[13]~3 .extended_lut = "off";
defparam \M_wr_data_unfiltered[13]~3 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \M_wr_data_unfiltered[13]~3 .shared_arith = "off";

dffeas \W_wr_data[13] (
	.clk(clk_clk),
	.d(\M_wr_data_unfiltered[13]~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\W_wr_data[13]~q ),
	.prn(vcc));
defparam \W_wr_data[13] .is_wysiwyg = "true";
defparam \W_wr_data[13] .power_up = "low";

cyclonev_lcell_comb \D_src1_prelim[13]~6 (
	.dataa(!\M_wr_data_unfiltered[13]~3_combout ),
	.datab(!\D_src1_hazard_M~combout ),
	.datac(!\D_src1_hazard_W~combout ),
	.datad(!\W_wr_data[13]~q ),
	.datae(!\processor_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[13] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_prelim[13]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src1_prelim[13]~6 .extended_lut = "off";
defparam \D_src1_prelim[13]~6 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \D_src1_prelim[13]~6 .shared_arith = "off";

dffeas \E_src1_prelim[13] (
	.clk(clk_clk),
	.d(\D_src1_prelim[13]~6_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_src1_prelim[13]~q ),
	.prn(vcc));
defparam \E_src1_prelim[13] .is_wysiwyg = "true";
defparam \E_src1_prelim[13] .power_up = "low";

cyclonev_lcell_comb \E_src1[13]~12 (
	.dataa(!\E_src1_hazard_M~q ),
	.datab(!\M_wr_data_unfiltered[13]~3_combout ),
	.datac(!\E_src1_prelim[13]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_src1[13]~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_src1[13]~12 .extended_lut = "off";
defparam \E_src1[13]~12 .lut_mask = 64'h2727272727272727;
defparam \E_src1[13]~12 .shared_arith = "off";

cyclonev_lcell_comb \M_shift_rot_result_nxt[13]~7 (
	.dataa(!\M_shift_rot_stall~q ),
	.datab(!\M_shift_rot_result[12]~q ),
	.datac(!\M_shift_rot_result[14]~q ),
	.datad(!\E_src1[13]~12_combout ),
	.datae(!\M_ctrl_shift_rot_right~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_shift_rot_result_nxt[13]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_shift_rot_result_nxt[13]~7 .extended_lut = "off";
defparam \M_shift_rot_result_nxt[13]~7 .lut_mask = 64'h7FFFBFFF7FFFBFFF;
defparam \M_shift_rot_result_nxt[13]~7 .shared_arith = "off";

dffeas \M_shift_rot_result[13] (
	.clk(clk_clk),
	.d(\M_shift_rot_result_nxt[13]~7_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\M_shift_rot_result[13]~q ),
	.prn(vcc));
defparam \M_shift_rot_result[13] .is_wysiwyg = "true";
defparam \M_shift_rot_result[13] .power_up = "low";

cyclonev_lcell_comb \M_shift_rot_result_nxt[14]~6 (
	.dataa(!\M_shift_rot_stall~q ),
	.datab(!\M_shift_rot_result[15]~q ),
	.datac(!\E_src1[14]~11_combout ),
	.datad(!\M_shift_rot_result[13]~q ),
	.datae(!\M_ctrl_shift_rot_right~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_shift_rot_result_nxt[14]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_shift_rot_result_nxt[14]~6 .extended_lut = "off";
defparam \M_shift_rot_result_nxt[14]~6 .lut_mask = 64'h7FFFBFFF7FFFBFFF;
defparam \M_shift_rot_result_nxt[14]~6 .shared_arith = "off";

dffeas \M_shift_rot_result[14] (
	.clk(clk_clk),
	.d(\M_shift_rot_result_nxt[14]~6_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\M_shift_rot_result[14]~q ),
	.prn(vcc));
defparam \M_shift_rot_result[14] .is_wysiwyg = "true";
defparam \M_shift_rot_result[14] .power_up = "low";

cyclonev_lcell_comb \M_shift_rot_result_nxt[15]~5 (
	.dataa(!\M_shift_rot_stall~q ),
	.datab(!\M_shift_rot_result[16]~q ),
	.datac(!\E_src1[15]~10_combout ),
	.datad(!\M_shift_rot_result[14]~q ),
	.datae(!\M_ctrl_shift_rot_right~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_shift_rot_result_nxt[15]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_shift_rot_result_nxt[15]~5 .extended_lut = "off";
defparam \M_shift_rot_result_nxt[15]~5 .lut_mask = 64'h7FFFBFFF7FFFBFFF;
defparam \M_shift_rot_result_nxt[15]~5 .shared_arith = "off";

dffeas \M_shift_rot_result[15] (
	.clk(clk_clk),
	.d(\M_shift_rot_result_nxt[15]~5_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\M_shift_rot_result[15]~q ),
	.prn(vcc));
defparam \M_shift_rot_result[15] .is_wysiwyg = "true";
defparam \M_shift_rot_result[15] .power_up = "low";

cyclonev_lcell_comb \M_shift_rot_result_nxt[16]~4 (
	.dataa(!\M_shift_rot_stall~q ),
	.datab(!\E_src1[16]~9_combout ),
	.datac(!\M_shift_rot_result[15]~q ),
	.datad(!\M_ctrl_shift_rot_right~q ),
	.datae(!\M_shift_rot_result[17]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_shift_rot_result_nxt[16]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_shift_rot_result_nxt[16]~4 .extended_lut = "off";
defparam \M_shift_rot_result_nxt[16]~4 .lut_mask = 64'h7FBFFFFF7FBFFFFF;
defparam \M_shift_rot_result_nxt[16]~4 .shared_arith = "off";

dffeas \M_shift_rot_result[16] (
	.clk(clk_clk),
	.d(\M_shift_rot_result_nxt[16]~4_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\M_shift_rot_result[16]~q ),
	.prn(vcc));
defparam \M_shift_rot_result[16] .is_wysiwyg = "true";
defparam \M_shift_rot_result[16] .power_up = "low";

dffeas \W_wr_data[17] (
	.clk(clk_clk),
	.d(\M_wr_data_unfiltered[17]~18_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\W_wr_data[17]~q ),
	.prn(vcc));
defparam \W_wr_data[17] .is_wysiwyg = "true";
defparam \W_wr_data[17] .power_up = "low";

cyclonev_lcell_comb \D_src1_prelim[17]~18 (
	.dataa(!\M_wr_data_unfiltered[17]~18_combout ),
	.datab(!\D_src1_hazard_M~combout ),
	.datac(!\D_src1_hazard_W~combout ),
	.datad(!\W_wr_data[17]~q ),
	.datae(!\processor_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[17] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_prelim[17]~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src1_prelim[17]~18 .extended_lut = "off";
defparam \D_src1_prelim[17]~18 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \D_src1_prelim[17]~18 .shared_arith = "off";

dffeas \E_src1_prelim[17] (
	.clk(clk_clk),
	.d(\D_src1_prelim[17]~18_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_src1_prelim[17]~q ),
	.prn(vcc));
defparam \E_src1_prelim[17] .is_wysiwyg = "true";
defparam \E_src1_prelim[17] .power_up = "low";

cyclonev_lcell_comb \E_src1[17]~32 (
	.dataa(!\E_src1_hazard_M~q ),
	.datab(!\M_wr_data_unfiltered[17]~18_combout ),
	.datac(!\E_src1_prelim[17]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_src1[17]~32_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_src1[17]~32 .extended_lut = "off";
defparam \E_src1[17]~32 .lut_mask = 64'h2727272727272727;
defparam \E_src1[17]~32 .shared_arith = "off";

cyclonev_lcell_comb \M_shift_rot_result_nxt[17]~18 (
	.dataa(!\M_shift_rot_stall~q ),
	.datab(!\M_shift_rot_result[16]~q ),
	.datac(!\M_ctrl_shift_rot_right~q ),
	.datad(!\M_shift_rot_result[18]~q ),
	.datae(!\E_src1[17]~32_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_shift_rot_result_nxt[17]~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_shift_rot_result_nxt[17]~18 .extended_lut = "off";
defparam \M_shift_rot_result_nxt[17]~18 .lut_mask = 64'h7BFFFFFF7BFFFFFF;
defparam \M_shift_rot_result_nxt[17]~18 .shared_arith = "off";

dffeas \M_shift_rot_result[17] (
	.clk(clk_clk),
	.d(\M_shift_rot_result_nxt[17]~18_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\M_shift_rot_result[17]~q ),
	.prn(vcc));
defparam \M_shift_rot_result[17] .is_wysiwyg = "true";
defparam \M_shift_rot_result[17] .power_up = "low";

dffeas \av_ld_data_aligned_or_div[17] (
	.clk(clk_clk),
	.d(\av_fill_bit~0_combout ),
	.asdata(\d_readdata_d1[17]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\M_iw[4]~q ),
	.ena(vcc),
	.q(\av_ld_data_aligned_or_div[17]~q ),
	.prn(vcc));
defparam \av_ld_data_aligned_or_div[17] .is_wysiwyg = "true";
defparam \av_ld_data_aligned_or_div[17] .power_up = "low";

cyclonev_lcell_comb \F_iw[7]~27 (
	.dataa(!\intr_req~0_combout ),
	.datab(!\processor_cpu_ic_data|the_altsyncram|auto_generated|q_b[7] ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[7]~27_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[7]~27 .extended_lut = "off";
defparam \F_iw[7]~27 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \F_iw[7]~27 .shared_arith = "off";

dffeas \D_iw[7] (
	.clk(clk_clk),
	.d(\F_iw[7]~27_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\F_iw~1_combout ),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\D_iw[7]~q ),
	.prn(vcc));
defparam \D_iw[7] .is_wysiwyg = "true";
defparam \D_iw[7] .power_up = "low";

dffeas \E_src2_imm[17] (
	.clk(clk_clk),
	.d(\D_iw[21]~q ),
	.asdata(\D_iw[7]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\D_ctrl_unsigned_lo_imm16~combout ),
	.sload(\Equal171~0_combout ),
	.ena(\W_stall~combout ),
	.q(\E_src2_imm[17]~q ),
	.prn(vcc));
defparam \E_src2_imm[17] .is_wysiwyg = "true";
defparam \E_src2_imm[17] .power_up = "low";

cyclonev_lcell_comb \E_stw_data[16]~0 (
	.dataa(!M_alu_result_16),
	.datab(!\E_src2_hazard_M~q ),
	.datac(!\M_ctrl_shift_rot~q ),
	.datad(!\av_ld_or_div_done~q ),
	.datae(!\M_shift_rot_result[16]~q ),
	.dataf(!\av_ld_data_aligned_or_div[16]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_stw_data[16]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_stw_data[16]~0 .extended_lut = "off";
defparam \E_stw_data[16]~0 .lut_mask = 64'h7FF7FFFFFFFFFFFF;
defparam \E_stw_data[16]~0 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_prelim[16]~4 (
	.dataa(!\M_wr_data_unfiltered[16]~13_combout ),
	.datab(!\D_src2_hazard_M~combout ),
	.datac(!\D_src2_hazard_W~combout ),
	.datad(!\W_wr_data[16]~q ),
	.datae(!\processor_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[16] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_prelim[16]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_prelim[16]~4 .extended_lut = "off";
defparam \D_src2_prelim[16]~4 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \D_src2_prelim[16]~4 .shared_arith = "off";

dffeas \E_src2_prelim[16] (
	.clk(clk_clk),
	.d(\D_src2_prelim[16]~4_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_src2_prelim[16]~q ),
	.prn(vcc));
defparam \E_src2_prelim[16] .is_wysiwyg = "true";
defparam \E_src2_prelim[16] .power_up = "low";

cyclonev_lcell_comb \E_stw_data[16]~1 (
	.dataa(!\E_src2_hazard_M~q ),
	.datab(!\E_src2_prelim[16]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_stw_data[16]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_stw_data[16]~1 .extended_lut = "off";
defparam \E_stw_data[16]~1 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \E_stw_data[16]~1 .shared_arith = "off";

cyclonev_lcell_comb \E_stw_data[16]~2 (
	.dataa(!\E_stw_data[16]~0_combout ),
	.datab(!\E_stw_data[16]~1_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_stw_data[16]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_stw_data[16]~2 .extended_lut = "off";
defparam \E_stw_data[16]~2 .lut_mask = 64'h7777777777777777;
defparam \E_stw_data[16]~2 .shared_arith = "off";

dffeas \E_src2_imm[16] (
	.clk(clk_clk),
	.d(\D_iw[21]~q ),
	.asdata(\D_iw[6]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\D_ctrl_unsigned_lo_imm16~combout ),
	.sload(\Equal171~0_combout ),
	.ena(\W_stall~combout ),
	.q(\E_src2_imm[16]~q ),
	.prn(vcc));
defparam \E_src2_imm[16] .is_wysiwyg = "true";
defparam \E_src2_imm[16] .power_up = "low";

cyclonev_lcell_comb \D_src2_prelim[15]~5 (
	.dataa(!\M_wr_data_unfiltered[15]~1_combout ),
	.datab(!\D_src2_hazard_M~combout ),
	.datac(!\D_src2_hazard_W~combout ),
	.datad(!\W_wr_data[15]~q ),
	.datae(!\processor_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[15] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_prelim[15]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_prelim[15]~5 .extended_lut = "off";
defparam \D_src2_prelim[15]~5 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \D_src2_prelim[15]~5 .shared_arith = "off";

dffeas \E_src2_prelim[15] (
	.clk(clk_clk),
	.d(\D_src2_prelim[15]~5_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_src2_prelim[15]~q ),
	.prn(vcc));
defparam \E_src2_prelim[15] .is_wysiwyg = "true";
defparam \E_src2_prelim[15] .power_up = "low";

cyclonev_lcell_comb \E_stw_data[15]~3 (
	.dataa(!\E_src2_hazard_M~q ),
	.datab(!\M_wr_data_unfiltered[15]~1_combout ),
	.datac(!\E_src2_prelim[15]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_stw_data[15]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_stw_data[15]~3 .extended_lut = "off";
defparam \E_stw_data[15]~3 .lut_mask = 64'h2727272727272727;
defparam \E_stw_data[15]~3 .shared_arith = "off";

dffeas \E_src2_imm[15] (
	.clk(clk_clk),
	.d(\D_iw[21]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\D_ctrl_hi_imm16~0_combout ),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_src2_imm[15]~q ),
	.prn(vcc));
defparam \E_src2_imm[15] .is_wysiwyg = "true";
defparam \E_src2_imm[15] .power_up = "low";

cyclonev_lcell_comb \D_src2_prelim[14]~6 (
	.dataa(!\M_wr_data_unfiltered[14]~2_combout ),
	.datab(!\D_src2_hazard_M~combout ),
	.datac(!\D_src2_hazard_W~combout ),
	.datad(!\W_wr_data[14]~q ),
	.datae(!\processor_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[14] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_prelim[14]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_prelim[14]~6 .extended_lut = "off";
defparam \D_src2_prelim[14]~6 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \D_src2_prelim[14]~6 .shared_arith = "off";

dffeas \E_src2_prelim[14] (
	.clk(clk_clk),
	.d(\D_src2_prelim[14]~6_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_src2_prelim[14]~q ),
	.prn(vcc));
defparam \E_src2_prelim[14] .is_wysiwyg = "true";
defparam \E_src2_prelim[14] .power_up = "low";

cyclonev_lcell_comb \E_stw_data[14]~4 (
	.dataa(!\E_src2_hazard_M~q ),
	.datab(!\M_wr_data_unfiltered[14]~2_combout ),
	.datac(!\E_src2_prelim[14]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_stw_data[14]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_stw_data[14]~4 .extended_lut = "off";
defparam \E_stw_data[14]~4 .lut_mask = 64'h2727272727272727;
defparam \E_stw_data[14]~4 .shared_arith = "off";

dffeas \E_src2_imm[14] (
	.clk(clk_clk),
	.d(\D_iw[20]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\D_ctrl_hi_imm16~0_combout ),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_src2_imm[14]~q ),
	.prn(vcc));
defparam \E_src2_imm[14] .is_wysiwyg = "true";
defparam \E_src2_imm[14] .power_up = "low";

cyclonev_lcell_comb \D_src2_prelim[13]~7 (
	.dataa(!\M_wr_data_unfiltered[13]~3_combout ),
	.datab(!\D_src2_hazard_M~combout ),
	.datac(!\D_src2_hazard_W~combout ),
	.datad(!\W_wr_data[13]~q ),
	.datae(!\processor_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[13] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_prelim[13]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_prelim[13]~7 .extended_lut = "off";
defparam \D_src2_prelim[13]~7 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \D_src2_prelim[13]~7 .shared_arith = "off";

dffeas \E_src2_prelim[13] (
	.clk(clk_clk),
	.d(\D_src2_prelim[13]~7_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_src2_prelim[13]~q ),
	.prn(vcc));
defparam \E_src2_prelim[13] .is_wysiwyg = "true";
defparam \E_src2_prelim[13] .power_up = "low";

cyclonev_lcell_comb \E_stw_data[13]~13 (
	.dataa(!\E_src2_hazard_M~q ),
	.datab(!\M_wr_data_unfiltered[13]~3_combout ),
	.datac(!\E_src2_prelim[13]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_stw_data[13]~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_stw_data[13]~13 .extended_lut = "off";
defparam \E_stw_data[13]~13 .lut_mask = 64'h2727272727272727;
defparam \E_stw_data[13]~13 .shared_arith = "off";

cyclonev_lcell_comb \F_iw[19]~29 (
	.dataa(!\F_iw~1_combout ),
	.datab(!\intr_req~0_combout ),
	.datac(!\processor_cpu_ic_data|the_altsyncram|auto_generated|q_b[19] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[19]~29_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[19]~29 .extended_lut = "off";
defparam \F_iw[19]~29 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \F_iw[19]~29 .shared_arith = "off";

dffeas \D_iw[19] (
	.clk(clk_clk),
	.d(\F_iw[19]~29_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\D_iw[19]~q ),
	.prn(vcc));
defparam \D_iw[19] .is_wysiwyg = "true";
defparam \D_iw[19] .power_up = "low";

dffeas \E_src2_imm[13] (
	.clk(clk_clk),
	.d(\D_iw[19]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\D_ctrl_hi_imm16~0_combout ),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_src2_imm[13]~q ),
	.prn(vcc));
defparam \E_src2_imm[13] .is_wysiwyg = "true";
defparam \E_src2_imm[13] .power_up = "low";

cyclonev_lcell_comb \D_src2_prelim[12]~8 (
	.dataa(!\M_wr_data_unfiltered[12]~4_combout ),
	.datab(!\D_src2_hazard_M~combout ),
	.datac(!\D_src2_hazard_W~combout ),
	.datad(!\W_wr_data[12]~q ),
	.datae(!\processor_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[12] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_prelim[12]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_prelim[12]~8 .extended_lut = "off";
defparam \D_src2_prelim[12]~8 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \D_src2_prelim[12]~8 .shared_arith = "off";

dffeas \E_src2_prelim[12] (
	.clk(clk_clk),
	.d(\D_src2_prelim[12]~8_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_src2_prelim[12]~q ),
	.prn(vcc));
defparam \E_src2_prelim[12] .is_wysiwyg = "true";
defparam \E_src2_prelim[12] .power_up = "low";

cyclonev_lcell_comb \E_stw_data[12]~5 (
	.dataa(!\E_src2_hazard_M~q ),
	.datab(!\M_wr_data_unfiltered[12]~4_combout ),
	.datac(!\E_src2_prelim[12]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_stw_data[12]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_stw_data[12]~5 .extended_lut = "off";
defparam \E_stw_data[12]~5 .lut_mask = 64'h2727272727272727;
defparam \E_stw_data[12]~5 .shared_arith = "off";

dffeas \E_src2_imm[12] (
	.clk(clk_clk),
	.d(\D_iw[18]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\D_ctrl_hi_imm16~0_combout ),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_src2_imm[12]~q ),
	.prn(vcc));
defparam \E_src2_imm[12] .is_wysiwyg = "true";
defparam \E_src2_imm[12] .power_up = "low";

cyclonev_lcell_comb \D_src2_prelim[11]~9 (
	.dataa(!\M_wr_data_unfiltered[11]~5_combout ),
	.datab(!\D_src2_hazard_M~combout ),
	.datac(!\D_src2_hazard_W~combout ),
	.datad(!\W_wr_data[11]~q ),
	.datae(!\processor_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[11] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_prelim[11]~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_prelim[11]~9 .extended_lut = "off";
defparam \D_src2_prelim[11]~9 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \D_src2_prelim[11]~9 .shared_arith = "off";

dffeas \E_src2_prelim[11] (
	.clk(clk_clk),
	.d(\D_src2_prelim[11]~9_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_src2_prelim[11]~q ),
	.prn(vcc));
defparam \E_src2_prelim[11] .is_wysiwyg = "true";
defparam \E_src2_prelim[11] .power_up = "low";

cyclonev_lcell_comb \E_stw_data[11]~14 (
	.dataa(!\E_src2_hazard_M~q ),
	.datab(!\M_wr_data_unfiltered[11]~5_combout ),
	.datac(!\E_src2_prelim[11]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_stw_data[11]~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_stw_data[11]~14 .extended_lut = "off";
defparam \E_stw_data[11]~14 .lut_mask = 64'h2727272727272727;
defparam \E_stw_data[11]~14 .shared_arith = "off";

dffeas \E_src2_imm[11] (
	.clk(clk_clk),
	.d(\D_iw[17]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\D_ctrl_hi_imm16~0_combout ),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_src2_imm[11]~q ),
	.prn(vcc));
defparam \E_src2_imm[11] .is_wysiwyg = "true";
defparam \E_src2_imm[11] .power_up = "low";

cyclonev_lcell_comb \E_stw_data[10]~6 (
	.dataa(!M_alu_result_10),
	.datab(!\E_src2_hazard_M~q ),
	.datac(!\M_ctrl_shift_rot~q ),
	.datad(!\av_ld_or_div_done~q ),
	.datae(!\M_shift_rot_result[10]~q ),
	.dataf(!\av_ld_data_aligned_or_div[10]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_stw_data[10]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_stw_data[10]~6 .extended_lut = "off";
defparam \E_stw_data[10]~6 .lut_mask = 64'h7FF7FFFFFFFFFFFF;
defparam \E_stw_data[10]~6 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_prelim[10]~10 (
	.dataa(!\M_wr_data_unfiltered[10]~14_combout ),
	.datab(!\D_src2_hazard_M~combout ),
	.datac(!\D_src2_hazard_W~combout ),
	.datad(!\W_wr_data[10]~q ),
	.datae(!\processor_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[10] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_prelim[10]~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_prelim[10]~10 .extended_lut = "off";
defparam \D_src2_prelim[10]~10 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \D_src2_prelim[10]~10 .shared_arith = "off";

dffeas \E_src2_prelim[10] (
	.clk(clk_clk),
	.d(\D_src2_prelim[10]~10_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_src2_prelim[10]~q ),
	.prn(vcc));
defparam \E_src2_prelim[10] .is_wysiwyg = "true";
defparam \E_src2_prelim[10] .power_up = "low";

cyclonev_lcell_comb \E_stw_data[10]~7 (
	.dataa(!\E_src2_hazard_M~q ),
	.datab(!\E_src2_prelim[10]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_stw_data[10]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_stw_data[10]~7 .extended_lut = "off";
defparam \E_stw_data[10]~7 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \E_stw_data[10]~7 .shared_arith = "off";

cyclonev_lcell_comb \E_stw_data[10]~8 (
	.dataa(!\E_stw_data[10]~6_combout ),
	.datab(!\E_stw_data[10]~7_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_stw_data[10]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_stw_data[10]~8 .extended_lut = "off";
defparam \E_stw_data[10]~8 .lut_mask = 64'h7777777777777777;
defparam \E_stw_data[10]~8 .shared_arith = "off";

dffeas \E_src2_imm[10] (
	.clk(clk_clk),
	.d(\D_iw[16]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\D_ctrl_hi_imm16~0_combout ),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_src2_imm[10]~q ),
	.prn(vcc));
defparam \E_src2_imm[10] .is_wysiwyg = "true";
defparam \E_src2_imm[10] .power_up = "low";

cyclonev_lcell_comb \D_src2_prelim[9]~11 (
	.dataa(!\M_wr_data_unfiltered[9]~6_combout ),
	.datab(!\D_src2_hazard_M~combout ),
	.datac(!\D_src2_hazard_W~combout ),
	.datad(!\W_wr_data[9]~q ),
	.datae(!\processor_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[9] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_prelim[9]~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_prelim[9]~11 .extended_lut = "off";
defparam \D_src2_prelim[9]~11 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \D_src2_prelim[9]~11 .shared_arith = "off";

dffeas \E_src2_prelim[9] (
	.clk(clk_clk),
	.d(\D_src2_prelim[9]~11_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_src2_prelim[9]~q ),
	.prn(vcc));
defparam \E_src2_prelim[9] .is_wysiwyg = "true";
defparam \E_src2_prelim[9] .power_up = "low";

cyclonev_lcell_comb \E_stw_data[9]~12 (
	.dataa(!\E_src2_hazard_M~q ),
	.datab(!\M_wr_data_unfiltered[9]~6_combout ),
	.datac(!\E_src2_prelim[9]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_stw_data[9]~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_stw_data[9]~12 .extended_lut = "off";
defparam \E_stw_data[9]~12 .lut_mask = 64'h2727272727272727;
defparam \E_stw_data[9]~12 .shared_arith = "off";

dffeas \E_src2_imm[9] (
	.clk(clk_clk),
	.d(\D_iw[15]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\D_ctrl_hi_imm16~0_combout ),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_src2_imm[9]~q ),
	.prn(vcc));
defparam \E_src2_imm[9] .is_wysiwyg = "true";
defparam \E_src2_imm[9] .power_up = "low";

cyclonev_lcell_comb \E_stw_data[8]~9 (
	.dataa(!M_alu_result_8),
	.datab(!\E_src2_hazard_M~q ),
	.datac(!\M_ctrl_shift_rot~q ),
	.datad(!\av_ld_or_div_done~q ),
	.datae(!\M_shift_rot_result[8]~q ),
	.dataf(!\av_ld_data_aligned_or_div[8]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_stw_data[8]~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_stw_data[8]~9 .extended_lut = "off";
defparam \E_stw_data[8]~9 .lut_mask = 64'h7FF7FFFFFFFFFFFF;
defparam \E_stw_data[8]~9 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_prelim[8]~12 (
	.dataa(!\M_wr_data_unfiltered[8]~15_combout ),
	.datab(!\D_src2_hazard_M~combout ),
	.datac(!\D_src2_hazard_W~combout ),
	.datad(!\W_wr_data[8]~q ),
	.datae(!\processor_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[8] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_prelim[8]~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_prelim[8]~12 .extended_lut = "off";
defparam \D_src2_prelim[8]~12 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \D_src2_prelim[8]~12 .shared_arith = "off";

dffeas \E_src2_prelim[8] (
	.clk(clk_clk),
	.d(\D_src2_prelim[8]~12_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_src2_prelim[8]~q ),
	.prn(vcc));
defparam \E_src2_prelim[8] .is_wysiwyg = "true";
defparam \E_src2_prelim[8] .power_up = "low";

cyclonev_lcell_comb \E_stw_data[8]~10 (
	.dataa(!\E_src2_hazard_M~q ),
	.datab(!\E_src2_prelim[8]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_stw_data[8]~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_stw_data[8]~10 .extended_lut = "off";
defparam \E_stw_data[8]~10 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \E_stw_data[8]~10 .shared_arith = "off";

cyclonev_lcell_comb \E_stw_data[8]~11 (
	.dataa(!\E_stw_data[8]~9_combout ),
	.datab(!\E_stw_data[8]~10_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_stw_data[8]~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_stw_data[8]~11 .extended_lut = "off";
defparam \E_stw_data[8]~11 .lut_mask = 64'h7777777777777777;
defparam \E_stw_data[8]~11 .shared_arith = "off";

dffeas \E_src2_imm[8] (
	.clk(clk_clk),
	.d(\D_iw[14]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\D_ctrl_hi_imm16~0_combout ),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_src2_imm[8]~q ),
	.prn(vcc));
defparam \E_src2_imm[8] .is_wysiwyg = "true";
defparam \E_src2_imm[8] .power_up = "low";

cyclonev_lcell_comb \D_src2_prelim[7]~13 (
	.dataa(!\M_wr_data_unfiltered[7]~7_combout ),
	.datab(!\D_src2_hazard_M~combout ),
	.datac(!\D_src2_hazard_W~combout ),
	.datad(!\W_wr_data[7]~q ),
	.datae(!\processor_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[7] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_prelim[7]~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_prelim[7]~13 .extended_lut = "off";
defparam \D_src2_prelim[7]~13 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \D_src2_prelim[7]~13 .shared_arith = "off";

dffeas \E_src2_prelim[7] (
	.clk(clk_clk),
	.d(\D_src2_prelim[7]~13_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_src2_prelim[7]~q ),
	.prn(vcc));
defparam \E_src2_prelim[7] .is_wysiwyg = "true";
defparam \E_src2_prelim[7] .power_up = "low";

cyclonev_lcell_comb \E_stb_data[7]~15 (
	.dataa(!\E_src2_hazard_M~q ),
	.datab(!\M_wr_data_unfiltered[7]~7_combout ),
	.datac(!\E_src2_prelim[7]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_stb_data[7]~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_stb_data[7]~15 .extended_lut = "off";
defparam \E_stb_data[7]~15 .lut_mask = 64'h2727272727272727;
defparam \E_stb_data[7]~15 .shared_arith = "off";

dffeas \E_src2_imm[7] (
	.clk(clk_clk),
	.d(\D_iw[13]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\D_ctrl_hi_imm16~0_combout ),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_src2_imm[7]~q ),
	.prn(vcc));
defparam \E_src2_imm[7] .is_wysiwyg = "true";
defparam \E_src2_imm[7] .power_up = "low";

cyclonev_lcell_comb \E_stb_data[6]~6 (
	.dataa(!M_alu_result_6),
	.datab(!\E_src2_hazard_M~q ),
	.datac(!\M_ctrl_shift_rot~q ),
	.datad(!\av_ld_or_div_done~q ),
	.datae(!\M_shift_rot_result[6]~q ),
	.dataf(!\av_ld_data_aligned_or_div[6]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_stb_data[6]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_stb_data[6]~6 .extended_lut = "off";
defparam \E_stb_data[6]~6 .lut_mask = 64'h7FF7FFFFFFFFFFFF;
defparam \E_stb_data[6]~6 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_prelim[6]~3 (
	.dataa(!\M_wr_data_unfiltered[6]~12_combout ),
	.datab(!\D_src2_hazard_M~combout ),
	.datac(!\D_src2_hazard_W~combout ),
	.datad(!\W_wr_data[6]~q ),
	.datae(!\processor_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[6] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_prelim[6]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_prelim[6]~3 .extended_lut = "off";
defparam \D_src2_prelim[6]~3 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \D_src2_prelim[6]~3 .shared_arith = "off";

dffeas \E_src2_prelim[6] (
	.clk(clk_clk),
	.d(\D_src2_prelim[6]~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_src2_prelim[6]~q ),
	.prn(vcc));
defparam \E_src2_prelim[6] .is_wysiwyg = "true";
defparam \E_src2_prelim[6] .power_up = "low";

cyclonev_lcell_comb \E_stb_data[6]~7 (
	.dataa(!\E_src2_hazard_M~q ),
	.datab(!\E_src2_prelim[6]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_stb_data[6]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_stb_data[6]~7 .extended_lut = "off";
defparam \E_stb_data[6]~7 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \E_stb_data[6]~7 .shared_arith = "off";

cyclonev_lcell_comb \E_stb_data[6]~8 (
	.dataa(!\E_stb_data[6]~6_combout ),
	.datab(!\E_stb_data[6]~7_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_stb_data[6]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_stb_data[6]~8 .extended_lut = "off";
defparam \E_stb_data[6]~8 .lut_mask = 64'h7777777777777777;
defparam \E_stb_data[6]~8 .shared_arith = "off";

dffeas \E_src2_imm[6] (
	.clk(clk_clk),
	.d(\D_iw[12]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\D_ctrl_hi_imm16~0_combout ),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_src2_imm[6]~q ),
	.prn(vcc));
defparam \E_src2_imm[6] .is_wysiwyg = "true";
defparam \E_src2_imm[6] .power_up = "low";

cyclonev_lcell_comb \D_src2_prelim[5]~1 (
	.dataa(!\M_wr_data_unfiltered[5]~0_combout ),
	.datab(!\D_src2_hazard_M~combout ),
	.datac(!\D_src2_hazard_W~combout ),
	.datad(!\W_wr_data[5]~q ),
	.datae(!\processor_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[5] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_prelim[5]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_prelim[5]~1 .extended_lut = "off";
defparam \D_src2_prelim[5]~1 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \D_src2_prelim[5]~1 .shared_arith = "off";

dffeas \E_src2_prelim[5] (
	.clk(clk_clk),
	.d(\D_src2_prelim[5]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_src2_prelim[5]~q ),
	.prn(vcc));
defparam \E_src2_prelim[5] .is_wysiwyg = "true";
defparam \E_src2_prelim[5] .power_up = "low";

cyclonev_lcell_comb \E_stb_data[5]~14 (
	.dataa(!\E_src2_hazard_M~q ),
	.datab(!\M_wr_data_unfiltered[5]~0_combout ),
	.datac(!\E_src2_prelim[5]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_stb_data[5]~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_stb_data[5]~14 .extended_lut = "off";
defparam \E_stb_data[5]~14 .lut_mask = 64'h2727272727272727;
defparam \E_stb_data[5]~14 .shared_arith = "off";

dffeas \E_src2_imm[5] (
	.clk(clk_clk),
	.d(\D_iw[11]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\D_ctrl_hi_imm16~0_combout ),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_src2_imm[5]~q ),
	.prn(vcc));
defparam \E_src2_imm[5] .is_wysiwyg = "true";
defparam \E_src2_imm[5] .power_up = "low";

cyclonev_lcell_comb \E_stb_data[4]~3 (
	.dataa(!M_alu_result_4),
	.datab(!\E_src2_hazard_M~q ),
	.datac(!\M_ctrl_shift_rot~q ),
	.datad(!\av_ld_or_div_done~q ),
	.datae(!\M_shift_rot_result[4]~q ),
	.dataf(!\av_ld_data_aligned_or_div[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_stb_data[4]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_stb_data[4]~3 .extended_lut = "off";
defparam \E_stb_data[4]~3 .lut_mask = 64'h7FF7FFFFFFFFFFFF;
defparam \E_stb_data[4]~3 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_prelim[4]~2 (
	.dataa(!\M_wr_data_unfiltered[4]~11_combout ),
	.datab(!\D_src2_hazard_M~combout ),
	.datac(!\D_src2_hazard_W~combout ),
	.datad(!\W_wr_data[4]~q ),
	.datae(!\processor_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[4] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_prelim[4]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_prelim[4]~2 .extended_lut = "off";
defparam \D_src2_prelim[4]~2 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \D_src2_prelim[4]~2 .shared_arith = "off";

dffeas \E_src2_prelim[4] (
	.clk(clk_clk),
	.d(\D_src2_prelim[4]~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_src2_prelim[4]~q ),
	.prn(vcc));
defparam \E_src2_prelim[4] .is_wysiwyg = "true";
defparam \E_src2_prelim[4] .power_up = "low";

cyclonev_lcell_comb \E_stb_data[4]~4 (
	.dataa(!\E_src2_hazard_M~q ),
	.datab(!\E_src2_prelim[4]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_stb_data[4]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_stb_data[4]~4 .extended_lut = "off";
defparam \E_stb_data[4]~4 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \E_stb_data[4]~4 .shared_arith = "off";

cyclonev_lcell_comb \E_stb_data[4]~5 (
	.dataa(!\E_stb_data[4]~3_combout ),
	.datab(!\E_stb_data[4]~4_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_stb_data[4]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_stb_data[4]~5 .extended_lut = "off";
defparam \E_stb_data[4]~5 .lut_mask = 64'h7777777777777777;
defparam \E_stb_data[4]~5 .shared_arith = "off";

dffeas \E_src2_imm[4] (
	.clk(clk_clk),
	.d(\D_iw[10]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\D_ctrl_hi_imm16~0_combout ),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_src2_imm[4]~q ),
	.prn(vcc));
defparam \E_src2_imm[4] .is_wysiwyg = "true";
defparam \E_src2_imm[4] .power_up = "low";

dffeas \W_wr_data[3] (
	.clk(clk_clk),
	.d(\M_wr_data_unfiltered[3]~8_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\W_wr_data[3]~q ),
	.prn(vcc));
defparam \W_wr_data[3] .is_wysiwyg = "true";
defparam \W_wr_data[3] .power_up = "low";

cyclonev_lcell_comb \D_src2_prelim[3]~14 (
	.dataa(!\M_wr_data_unfiltered[3]~8_combout ),
	.datab(!\D_src2_hazard_M~combout ),
	.datac(!\D_src2_hazard_W~combout ),
	.datad(!\W_wr_data[3]~q ),
	.datae(!\processor_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[3] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_prelim[3]~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_prelim[3]~14 .extended_lut = "off";
defparam \D_src2_prelim[3]~14 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \D_src2_prelim[3]~14 .shared_arith = "off";

dffeas \E_src2_prelim[3] (
	.clk(clk_clk),
	.d(\D_src2_prelim[3]~14_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_src2_prelim[3]~q ),
	.prn(vcc));
defparam \E_src2_prelim[3] .is_wysiwyg = "true";
defparam \E_src2_prelim[3] .power_up = "low";

cyclonev_lcell_comb \E_stb_data[3]~13 (
	.dataa(!\E_src2_hazard_M~q ),
	.datab(!\M_wr_data_unfiltered[3]~8_combout ),
	.datac(!\E_src2_prelim[3]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_stb_data[3]~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_stb_data[3]~13 .extended_lut = "off";
defparam \E_stb_data[3]~13 .lut_mask = 64'h2727272727272727;
defparam \E_stb_data[3]~13 .shared_arith = "off";

cyclonev_lcell_comb \F_iw[9]~32 (
	.dataa(!\intr_req~0_combout ),
	.datab(!\processor_cpu_ic_data|the_altsyncram|auto_generated|q_b[9] ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[9]~32_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[9]~32 .extended_lut = "off";
defparam \F_iw[9]~32 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \F_iw[9]~32 .shared_arith = "off";

dffeas \D_iw[9] (
	.clk(clk_clk),
	.d(\F_iw[9]~32_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\F_iw~1_combout ),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\D_iw[9]~q ),
	.prn(vcc));
defparam \D_iw[9] .is_wysiwyg = "true";
defparam \D_iw[9] .power_up = "low";

dffeas \E_src2_imm[3] (
	.clk(clk_clk),
	.d(\D_iw[9]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\D_ctrl_hi_imm16~0_combout ),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_src2_imm[3]~q ),
	.prn(vcc));
defparam \E_src2_imm[3] .is_wysiwyg = "true";
defparam \E_src2_imm[3] .power_up = "low";

dffeas \d_readdata_d1[2] (
	.clk(clk_clk),
	.d(d_readdata[2]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d_readdata_d1[2]~q ),
	.prn(vcc));
defparam \d_readdata_d1[2] .is_wysiwyg = "true";
defparam \d_readdata_d1[2] .power_up = "low";

cyclonev_lcell_comb \av_ld_byte0_data[2]~6 (
	.dataa(!\d_readdata_d1[2]~q ),
	.datab(!\d_readdata_d1[18]~q ),
	.datac(!\d_readdata_d1[10]~q ),
	.datad(!\d_readdata_d1[26]~q ),
	.datae(!\M_ld_align_sh16~combout ),
	.dataf(!\M_ld_align_sh8~combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_ld_byte0_data[2]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_ld_byte0_data[2]~6 .extended_lut = "off";
defparam \av_ld_byte0_data[2]~6 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \av_ld_byte0_data[2]~6 .shared_arith = "off";

dffeas \av_ld_data_aligned_or_div[2] (
	.clk(clk_clk),
	.d(\av_ld_byte0_data[2]~6_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\av_ld_data_aligned_or_div[2]~q ),
	.prn(vcc));
defparam \av_ld_data_aligned_or_div[2] .is_wysiwyg = "true";
defparam \av_ld_data_aligned_or_div[2] .power_up = "low";

cyclonev_lcell_comb \E_stb_data[2]~9 (
	.dataa(!M_alu_result_2),
	.datab(!\E_src2_hazard_M~q ),
	.datac(!\M_ctrl_shift_rot~q ),
	.datad(!\av_ld_or_div_done~q ),
	.datae(!\M_shift_rot_result[2]~q ),
	.dataf(!\av_ld_data_aligned_or_div[2]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_stb_data[2]~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_stb_data[2]~9 .extended_lut = "off";
defparam \E_stb_data[2]~9 .lut_mask = 64'h7FF7FFFFFFFFFFFF;
defparam \E_stb_data[2]~9 .shared_arith = "off";

cyclonev_lcell_comb \M_wr_data_unfiltered[2]~16 (
	.dataa(!M_alu_result_2),
	.datab(!\M_ctrl_shift_rot~q ),
	.datac(!\av_ld_or_div_done~q ),
	.datad(!\M_shift_rot_result[2]~q ),
	.datae(!\av_ld_data_aligned_or_div[2]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_wr_data_unfiltered[2]~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_wr_data_unfiltered[2]~16 .extended_lut = "off";
defparam \M_wr_data_unfiltered[2]~16 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \M_wr_data_unfiltered[2]~16 .shared_arith = "off";

dffeas \W_wr_data[2] (
	.clk(clk_clk),
	.d(\M_wr_data_unfiltered[2]~16_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\W_wr_data[2]~q ),
	.prn(vcc));
defparam \W_wr_data[2] .is_wysiwyg = "true";
defparam \W_wr_data[2] .power_up = "low";

cyclonev_lcell_comb \D_src2_prelim[2]~15 (
	.dataa(!\M_wr_data_unfiltered[2]~16_combout ),
	.datab(!\D_src2_hazard_M~combout ),
	.datac(!\D_src2_hazard_W~combout ),
	.datad(!\W_wr_data[2]~q ),
	.datae(!\processor_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[2] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_prelim[2]~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_prelim[2]~15 .extended_lut = "off";
defparam \D_src2_prelim[2]~15 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \D_src2_prelim[2]~15 .shared_arith = "off";

dffeas \E_src2_prelim[2] (
	.clk(clk_clk),
	.d(\D_src2_prelim[2]~15_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_src2_prelim[2]~q ),
	.prn(vcc));
defparam \E_src2_prelim[2] .is_wysiwyg = "true";
defparam \E_src2_prelim[2] .power_up = "low";

cyclonev_lcell_comb \E_stb_data[2]~10 (
	.dataa(!\E_src2_hazard_M~q ),
	.datab(!\E_src2_prelim[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_stb_data[2]~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_stb_data[2]~10 .extended_lut = "off";
defparam \E_stb_data[2]~10 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \E_stb_data[2]~10 .shared_arith = "off";

cyclonev_lcell_comb \E_stb_data[2]~11 (
	.dataa(!\E_stb_data[2]~9_combout ),
	.datab(!\E_stb_data[2]~10_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_stb_data[2]~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_stb_data[2]~11 .extended_lut = "off";
defparam \E_stb_data[2]~11 .lut_mask = 64'h7777777777777777;
defparam \E_stb_data[2]~11 .shared_arith = "off";

dffeas \E_src2_imm[2] (
	.clk(clk_clk),
	.d(\D_iw[8]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\D_ctrl_hi_imm16~0_combout ),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_src2_imm[2]~q ),
	.prn(vcc));
defparam \E_src2_imm[2] .is_wysiwyg = "true";
defparam \E_src2_imm[2] .power_up = "low";

cyclonev_lcell_comb \E_src1[2]~24 (
	.dataa(!M_alu_result_2),
	.datab(!\M_ctrl_shift_rot~q ),
	.datac(!\av_ld_or_div_done~q ),
	.datad(!\E_src1_hazard_M~q ),
	.datae(!\M_shift_rot_result[2]~q ),
	.dataf(!\av_ld_data_aligned_or_div[2]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_src1[2]~24_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_src1[2]~24 .extended_lut = "off";
defparam \E_src1[2]~24 .lut_mask = 64'h7DFFFFFFFFFFFFFF;
defparam \E_src1[2]~24 .shared_arith = "off";

cyclonev_lcell_comb \D_src1_prelim[2]~14 (
	.dataa(!\M_wr_data_unfiltered[2]~16_combout ),
	.datab(!\D_src1_hazard_M~combout ),
	.datac(!\D_src1_hazard_W~combout ),
	.datad(!\W_wr_data[2]~q ),
	.datae(!\processor_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[2] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_prelim[2]~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src1_prelim[2]~14 .extended_lut = "off";
defparam \D_src1_prelim[2]~14 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \D_src1_prelim[2]~14 .shared_arith = "off";

dffeas \E_src1_prelim[2] (
	.clk(clk_clk),
	.d(\D_src1_prelim[2]~14_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_src1_prelim[2]~q ),
	.prn(vcc));
defparam \E_src1_prelim[2] .is_wysiwyg = "true";
defparam \E_src1_prelim[2] .power_up = "low";

cyclonev_lcell_comb \E_src1[2]~25 (
	.dataa(!\E_src1_hazard_M~q ),
	.datab(!\E_src1_prelim[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_src1[2]~25_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_src1[2]~25 .extended_lut = "off";
defparam \E_src1[2]~25 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \E_src1[2]~25 .shared_arith = "off";

cyclonev_lcell_comb \E_src1[2]~26 (
	.dataa(!\E_src1[2]~24_combout ),
	.datab(!\E_src1[2]~25_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_src1[2]~26_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_src1[2]~26 .extended_lut = "off";
defparam \E_src1[2]~26 .lut_mask = 64'h7777777777777777;
defparam \E_src1[2]~26 .shared_arith = "off";

dffeas \E_src2_imm[1] (
	.clk(clk_clk),
	.d(\D_iw[7]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\D_ctrl_hi_imm16~0_combout ),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_src2_imm[1]~q ),
	.prn(vcc));
defparam \E_src2_imm[1] .is_wysiwyg = "true";
defparam \E_src2_imm[1] .power_up = "low";

dffeas \W_wr_data[1] (
	.clk(clk_clk),
	.d(\M_wr_data_unfiltered[1]~9_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\W_wr_data[1]~q ),
	.prn(vcc));
defparam \W_wr_data[1] .is_wysiwyg = "true";
defparam \W_wr_data[1] .power_up = "low";

cyclonev_lcell_comb \D_src1_prelim[1]~16 (
	.dataa(!\M_wr_data_unfiltered[1]~9_combout ),
	.datab(!\D_src1_hazard_M~combout ),
	.datac(!\D_src1_hazard_W~combout ),
	.datad(!\W_wr_data[1]~q ),
	.datae(!\processor_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[1] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_prelim[1]~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src1_prelim[1]~16 .extended_lut = "off";
defparam \D_src1_prelim[1]~16 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \D_src1_prelim[1]~16 .shared_arith = "off";

dffeas \E_src1_prelim[1] (
	.clk(clk_clk),
	.d(\D_src1_prelim[1]~16_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_src1_prelim[1]~q ),
	.prn(vcc));
defparam \E_src1_prelim[1] .is_wysiwyg = "true";
defparam \E_src1_prelim[1] .power_up = "low";

cyclonev_lcell_comb \E_src1[1]~30 (
	.dataa(!\E_src1_hazard_M~q ),
	.datab(!\M_wr_data_unfiltered[1]~9_combout ),
	.datac(!\E_src1_prelim[1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_src1[1]~30_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_src1[1]~30 .extended_lut = "off";
defparam \E_src1[1]~30 .lut_mask = 64'h2727272727272727;
defparam \E_src1[1]~30 .shared_arith = "off";

dffeas \d_readdata_d1[0] (
	.clk(clk_clk),
	.d(d_readdata[0]),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d_readdata_d1[0]~q ),
	.prn(vcc));
defparam \d_readdata_d1[0] .is_wysiwyg = "true";
defparam \d_readdata_d1[0] .power_up = "low";

cyclonev_lcell_comb \av_ld_byte0_data[0]~0 (
	.dataa(!\d_readdata_d1[0]~q ),
	.datab(!\d_readdata_d1[16]~q ),
	.datac(!\d_readdata_d1[8]~q ),
	.datad(!\d_readdata_d1[24]~q ),
	.datae(!\M_ld_align_sh16~combout ),
	.dataf(!\M_ld_align_sh8~combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_ld_byte0_data[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_ld_byte0_data[0]~0 .extended_lut = "off";
defparam \av_ld_byte0_data[0]~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \av_ld_byte0_data[0]~0 .shared_arith = "off";

dffeas \av_ld_data_aligned_or_div[0] (
	.clk(clk_clk),
	.d(\av_ld_byte0_data[0]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\av_ld_data_aligned_or_div[0]~q ),
	.prn(vcc));
defparam \av_ld_data_aligned_or_div[0] .is_wysiwyg = "true";
defparam \av_ld_data_aligned_or_div[0] .power_up = "low";

cyclonev_lcell_comb \E_src1[0]~27 (
	.dataa(!\M_shift_rot_result[0]~q ),
	.datab(!\M_ctrl_shift_rot~q ),
	.datac(!\av_ld_data_aligned_or_div[0]~q ),
	.datad(!\av_ld_or_div_done~q ),
	.datae(!\M_alu_result[0]~q ),
	.dataf(!\E_src1_hazard_M~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_src1[0]~27_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_src1[0]~27 .extended_lut = "off";
defparam \E_src1[0]~27 .lut_mask = 64'h7FDFFFFFFFFFFFFF;
defparam \E_src1[0]~27 .shared_arith = "off";

dffeas \W_wr_data[0] (
	.clk(clk_clk),
	.d(\M_wr_data_unfiltered[0]~10_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\W_wr_data[0]~q ),
	.prn(vcc));
defparam \W_wr_data[0] .is_wysiwyg = "true";
defparam \W_wr_data[0] .power_up = "low";

cyclonev_lcell_comb \D_src1_prelim[0]~15 (
	.dataa(!\M_wr_data_unfiltered[0]~10_combout ),
	.datab(!\W_wr_data[0]~q ),
	.datac(!\D_src1_hazard_M~combout ),
	.datad(!\D_src1_hazard_W~combout ),
	.datae(!\processor_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[0] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_prelim[0]~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src1_prelim[0]~15 .extended_lut = "off";
defparam \D_src1_prelim[0]~15 .lut_mask = 64'h7FF7FFFF7FF7FFFF;
defparam \D_src1_prelim[0]~15 .shared_arith = "off";

dffeas \E_src1_prelim[0] (
	.clk(clk_clk),
	.d(\D_src1_prelim[0]~15_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_src1_prelim[0]~q ),
	.prn(vcc));
defparam \E_src1_prelim[0] .is_wysiwyg = "true";
defparam \E_src1_prelim[0] .power_up = "low";

cyclonev_lcell_comb \E_src1[0]~28 (
	.dataa(!\E_src1_hazard_M~q ),
	.datab(!\E_src1_prelim[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_src1[0]~28_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_src1[0]~28 .extended_lut = "off";
defparam \E_src1[0]~28 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \E_src1[0]~28 .shared_arith = "off";

cyclonev_lcell_comb \E_src1[0]~29 (
	.dataa(!\E_src1[0]~27_combout ),
	.datab(!\E_src1[0]~28_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_src1[0]~29_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_src1[0]~29 .extended_lut = "off";
defparam \E_src1[0]~29 .lut_mask = 64'h7777777777777777;
defparam \E_src1[0]~29 .shared_arith = "off";

cyclonev_lcell_comb \Add8~78 (
	.dataa(!\E_ctrl_alu_subtract~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\Add8~78_cout ),
	.shareout());
defparam \Add8~78 .extended_lut = "off";
defparam \Add8~78 .lut_mask = 64'h0000000000005555;
defparam \Add8~78 .shared_arith = "off";

cyclonev_lcell_comb \Add8~65 (
	.dataa(!\E_ctrl_alu_subtract~q ),
	.datab(!\E_ctrl_src2_choose_imm~q ),
	.datac(!\E_stb_data[0]~2_combout ),
	.datad(!\E_src2_imm[0]~q ),
	.datae(gnd),
	.dataf(!\E_src1[0]~29_combout ),
	.datag(gnd),
	.cin(\Add8~78_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add8~65_sumout ),
	.cout(\Add8~66 ),
	.shareout());
defparam \Add8~65 .extended_lut = "off";
defparam \Add8~65 .lut_mask = 64'h0000FF0000006996;
defparam \Add8~65 .shared_arith = "off";

cyclonev_lcell_comb \Add8~69 (
	.dataa(!\E_ctrl_alu_subtract~q ),
	.datab(!\E_ctrl_src2_choose_imm~q ),
	.datac(!\E_stb_data[1]~12_combout ),
	.datad(!\E_src2_imm[1]~q ),
	.datae(gnd),
	.dataf(!\E_src1[1]~30_combout ),
	.datag(gnd),
	.cin(\Add8~66 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add8~69_sumout ),
	.cout(\Add8~70 ),
	.shareout());
defparam \Add8~69 .extended_lut = "off";
defparam \Add8~69 .lut_mask = 64'h0000FF0000006996;
defparam \Add8~69 .shared_arith = "off";

cyclonev_lcell_comb \Add8~57 (
	.dataa(!\E_ctrl_alu_subtract~q ),
	.datab(!\E_ctrl_src2_choose_imm~q ),
	.datac(!\E_stb_data[2]~11_combout ),
	.datad(!\E_src2_imm[2]~q ),
	.datae(gnd),
	.dataf(!\E_src1[2]~26_combout ),
	.datag(gnd),
	.cin(\Add8~70 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add8~57_sumout ),
	.cout(\Add8~58 ),
	.shareout());
defparam \Add8~57 .extended_lut = "off";
defparam \Add8~57 .lut_mask = 64'h0000FF0000006996;
defparam \Add8~57 .shared_arith = "off";

cyclonev_lcell_comb \Add8~53 (
	.dataa(!\E_ctrl_alu_subtract~q ),
	.datab(!\E_ctrl_src2_choose_imm~q ),
	.datac(!\E_stb_data[3]~13_combout ),
	.datad(!\E_src2_imm[3]~q ),
	.datae(gnd),
	.dataf(!\E_src1[3]~23_combout ),
	.datag(gnd),
	.cin(\Add8~58 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add8~53_sumout ),
	.cout(\Add8~54 ),
	.shareout());
defparam \Add8~53 .extended_lut = "off";
defparam \Add8~53 .lut_mask = 64'h0000FF0000006996;
defparam \Add8~53 .shared_arith = "off";

cyclonev_lcell_comb \Add8~5 (
	.dataa(!\E_ctrl_alu_subtract~q ),
	.datab(!\E_ctrl_src2_choose_imm~q ),
	.datac(!\E_stb_data[4]~5_combout ),
	.datad(!\E_src2_imm[4]~q ),
	.datae(gnd),
	.dataf(!\E_src1[4]~3_combout ),
	.datag(gnd),
	.cin(\Add8~54 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add8~5_sumout ),
	.cout(\Add8~6 ),
	.shareout());
defparam \Add8~5 .extended_lut = "off";
defparam \Add8~5 .lut_mask = 64'h0000FF0000006996;
defparam \Add8~5 .shared_arith = "off";

cyclonev_lcell_comb \Add8~1 (
	.dataa(!\E_ctrl_alu_subtract~q ),
	.datab(!\E_ctrl_src2_choose_imm~q ),
	.datac(!\E_stb_data[5]~14_combout ),
	.datad(!\E_src2_imm[5]~q ),
	.datae(gnd),
	.dataf(!\E_src1[5]~0_combout ),
	.datag(gnd),
	.cin(\Add8~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add8~1_sumout ),
	.cout(\Add8~2 ),
	.shareout());
defparam \Add8~1 .extended_lut = "off";
defparam \Add8~1 .lut_mask = 64'h0000FF0000006996;
defparam \Add8~1 .shared_arith = "off";

cyclonev_lcell_comb \Add8~9 (
	.dataa(!\E_ctrl_alu_subtract~q ),
	.datab(!\E_ctrl_src2_choose_imm~q ),
	.datac(!\E_stb_data[6]~8_combout ),
	.datad(!\E_src2_imm[6]~q ),
	.datae(gnd),
	.dataf(!\E_src1[6]~6_combout ),
	.datag(gnd),
	.cin(\Add8~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add8~9_sumout ),
	.cout(\Add8~10 ),
	.shareout());
defparam \Add8~9 .extended_lut = "off";
defparam \Add8~9 .lut_mask = 64'h0000FF0000006996;
defparam \Add8~9 .shared_arith = "off";

cyclonev_lcell_comb \Add8~49 (
	.dataa(!\E_ctrl_alu_subtract~q ),
	.datab(!\E_ctrl_src2_choose_imm~q ),
	.datac(!\E_stb_data[7]~15_combout ),
	.datad(!\E_src2_imm[7]~q ),
	.datae(gnd),
	.dataf(!\E_src1[7]~22_combout ),
	.datag(gnd),
	.cin(\Add8~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add8~49_sumout ),
	.cout(\Add8~50 ),
	.shareout());
defparam \Add8~49 .extended_lut = "off";
defparam \Add8~49 .lut_mask = 64'h0000FF0000006996;
defparam \Add8~49 .shared_arith = "off";

cyclonev_lcell_comb \Add8~45 (
	.dataa(!\E_ctrl_alu_subtract~q ),
	.datab(!\E_ctrl_src2_choose_imm~q ),
	.datac(!\E_stw_data[8]~11_combout ),
	.datad(!\E_src2_imm[8]~q ),
	.datae(gnd),
	.dataf(!\E_src1[8]~21_combout ),
	.datag(gnd),
	.cin(\Add8~50 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add8~45_sumout ),
	.cout(\Add8~46 ),
	.shareout());
defparam \Add8~45 .extended_lut = "off";
defparam \Add8~45 .lut_mask = 64'h0000FF0000006996;
defparam \Add8~45 .shared_arith = "off";

cyclonev_lcell_comb \Add8~41 (
	.dataa(!\E_ctrl_alu_subtract~q ),
	.datab(!\E_ctrl_src2_choose_imm~q ),
	.datac(!\E_stw_data[9]~12_combout ),
	.datad(!\E_src2_imm[9]~q ),
	.datae(gnd),
	.dataf(!\E_src1[9]~18_combout ),
	.datag(gnd),
	.cin(\Add8~46 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add8~41_sumout ),
	.cout(\Add8~42 ),
	.shareout());
defparam \Add8~41 .extended_lut = "off";
defparam \Add8~41 .lut_mask = 64'h0000FF0000006996;
defparam \Add8~41 .shared_arith = "off";

cyclonev_lcell_comb \Add8~37 (
	.dataa(!\E_ctrl_alu_subtract~q ),
	.datab(!\E_ctrl_src2_choose_imm~q ),
	.datac(!\E_stw_data[10]~8_combout ),
	.datad(!\E_src2_imm[10]~q ),
	.datae(gnd),
	.dataf(!\E_src1[10]~17_combout ),
	.datag(gnd),
	.cin(\Add8~42 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add8~37_sumout ),
	.cout(\Add8~38 ),
	.shareout());
defparam \Add8~37 .extended_lut = "off";
defparam \Add8~37 .lut_mask = 64'h0000FF0000006996;
defparam \Add8~37 .shared_arith = "off";

cyclonev_lcell_comb \Add8~33 (
	.dataa(!\E_ctrl_alu_subtract~q ),
	.datab(!\E_ctrl_src2_choose_imm~q ),
	.datac(!\E_stw_data[11]~14_combout ),
	.datad(!\E_src2_imm[11]~q ),
	.datae(gnd),
	.dataf(!\E_src1[11]~14_combout ),
	.datag(gnd),
	.cin(\Add8~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add8~33_sumout ),
	.cout(\Add8~34 ),
	.shareout());
defparam \Add8~33 .extended_lut = "off";
defparam \Add8~33 .lut_mask = 64'h0000FF0000006996;
defparam \Add8~33 .shared_arith = "off";

cyclonev_lcell_comb \Add8~29 (
	.dataa(!\E_ctrl_alu_subtract~q ),
	.datab(!\E_ctrl_src2_choose_imm~q ),
	.datac(!\E_stw_data[12]~5_combout ),
	.datad(!\E_src2_imm[12]~q ),
	.datae(gnd),
	.dataf(!\E_src1[12]~13_combout ),
	.datag(gnd),
	.cin(\Add8~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add8~29_sumout ),
	.cout(\Add8~30 ),
	.shareout());
defparam \Add8~29 .extended_lut = "off";
defparam \Add8~29 .lut_mask = 64'h0000FF0000006996;
defparam \Add8~29 .shared_arith = "off";

cyclonev_lcell_comb \Add8~25 (
	.dataa(!\E_ctrl_alu_subtract~q ),
	.datab(!\E_ctrl_src2_choose_imm~q ),
	.datac(!\E_stw_data[13]~13_combout ),
	.datad(!\E_src2_imm[13]~q ),
	.datae(gnd),
	.dataf(!\E_src1[13]~12_combout ),
	.datag(gnd),
	.cin(\Add8~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add8~25_sumout ),
	.cout(\Add8~26 ),
	.shareout());
defparam \Add8~25 .extended_lut = "off";
defparam \Add8~25 .lut_mask = 64'h0000FF0000006996;
defparam \Add8~25 .shared_arith = "off";

cyclonev_lcell_comb \Add8~21 (
	.dataa(!\E_ctrl_alu_subtract~q ),
	.datab(!\E_ctrl_src2_choose_imm~q ),
	.datac(!\E_stw_data[14]~4_combout ),
	.datad(!\E_src2_imm[14]~q ),
	.datae(gnd),
	.dataf(!\E_src1[14]~11_combout ),
	.datag(gnd),
	.cin(\Add8~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add8~21_sumout ),
	.cout(\Add8~22 ),
	.shareout());
defparam \Add8~21 .extended_lut = "off";
defparam \Add8~21 .lut_mask = 64'h0000FF0000006996;
defparam \Add8~21 .shared_arith = "off";

cyclonev_lcell_comb \Add8~17 (
	.dataa(!\E_ctrl_alu_subtract~q ),
	.datab(!\E_ctrl_src2_choose_imm~q ),
	.datac(!\E_stw_data[15]~3_combout ),
	.datad(!\E_src2_imm[15]~q ),
	.datae(gnd),
	.dataf(!\E_src1[15]~10_combout ),
	.datag(gnd),
	.cin(\Add8~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add8~17_sumout ),
	.cout(\Add8~18 ),
	.shareout());
defparam \Add8~17 .extended_lut = "off";
defparam \Add8~17 .lut_mask = 64'h0000FF0000006996;
defparam \Add8~17 .shared_arith = "off";

cyclonev_lcell_comb \Add8~13 (
	.dataa(!\E_ctrl_alu_subtract~q ),
	.datab(!\E_ctrl_src2_choose_imm~q ),
	.datac(!\E_stw_data[16]~2_combout ),
	.datad(!\E_src2_imm[16]~q ),
	.datae(gnd),
	.dataf(!\E_src1[16]~9_combout ),
	.datag(gnd),
	.cin(\Add8~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add8~13_sumout ),
	.cout(\Add8~14 ),
	.shareout());
defparam \Add8~13 .extended_lut = "off";
defparam \Add8~13 .lut_mask = 64'h0000FF0000006996;
defparam \Add8~13 .shared_arith = "off";

cyclonev_lcell_comb \Add8~85 (
	.dataa(!\E_ctrl_alu_subtract~q ),
	.datab(!\E_ctrl_src2_choose_imm~q ),
	.datac(!\E_stw_data[17]~35_combout ),
	.datad(!\E_src2_imm[17]~q ),
	.datae(gnd),
	.dataf(!\E_src1[17]~32_combout ),
	.datag(gnd),
	.cin(\Add8~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add8~85_sumout ),
	.cout(\Add8~86 ),
	.shareout());
defparam \Add8~85 .extended_lut = "off";
defparam \Add8~85 .lut_mask = 64'h0000FF0000006996;
defparam \Add8~85 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_prelim[17]~18 (
	.dataa(!\M_wr_data_unfiltered[17]~18_combout ),
	.datab(!\D_src2_hazard_M~combout ),
	.datac(!\D_src2_hazard_W~combout ),
	.datad(!\W_wr_data[17]~q ),
	.datae(!\processor_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[17] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_prelim[17]~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_prelim[17]~18 .extended_lut = "off";
defparam \D_src2_prelim[17]~18 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \D_src2_prelim[17]~18 .shared_arith = "off";

dffeas \E_src2_prelim[17] (
	.clk(clk_clk),
	.d(\D_src2_prelim[17]~18_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_src2_prelim[17]~q ),
	.prn(vcc));
defparam \E_src2_prelim[17] .is_wysiwyg = "true";
defparam \E_src2_prelim[17] .power_up = "low";

cyclonev_lcell_comb \E_arith_src2[17]~13 (
	.dataa(!\E_src2_hazard_M~q ),
	.datab(!\E_ctrl_src2_choose_imm~q ),
	.datac(!\M_wr_data_unfiltered[17]~18_combout ),
	.datad(!\E_src2_imm[17]~q ),
	.datae(!\E_src2_prelim[17]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_arith_src2[17]~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_arith_src2[17]~13 .extended_lut = "off";
defparam \E_arith_src2[17]~13 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \E_arith_src2[17]~13 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[17]~28 (
	.dataa(!\E_compare_op[1]~q ),
	.datab(!\E_compare_op[0]~q ),
	.datac(!\E_arith_src2[17]~13_combout ),
	.datad(!\E_src1[17]~32_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[17]~28_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[17]~28 .extended_lut = "off";
defparam \E_alu_result[17]~28 .lut_mask = 64'h6996699669966996;
defparam \E_alu_result[17]~28 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[17]~29 (
	.dataa(!\E_ctrl_logic~q ),
	.datab(!\E_alu_result~0_combout ),
	.datac(!\Add8~85_sumout ),
	.datad(!\E_alu_result[17]~28_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[17]~29_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[17]~29 .extended_lut = "off";
defparam \E_alu_result[17]~29 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \E_alu_result[17]~29 .shared_arith = "off";

dffeas \M_alu_result[17] (
	.clk(clk_clk),
	.d(\E_alu_result[17]~29_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\M_alu_result[17]~q ),
	.prn(vcc));
defparam \M_alu_result[17] .is_wysiwyg = "true";
defparam \M_alu_result[17] .power_up = "low";

cyclonev_lcell_comb \M_wr_data_unfiltered[17]~18 (
	.dataa(!\M_ctrl_shift_rot~q ),
	.datab(!\av_ld_or_div_done~q ),
	.datac(!\M_shift_rot_result[17]~q ),
	.datad(!\av_ld_data_aligned_or_div[17]~q ),
	.datae(!\M_alu_result[17]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_wr_data_unfiltered[17]~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_wr_data_unfiltered[17]~18 .extended_lut = "off";
defparam \M_wr_data_unfiltered[17]~18 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \M_wr_data_unfiltered[17]~18 .shared_arith = "off";

cyclonev_lcell_comb \E_stw_data[17]~35 (
	.dataa(!\E_src2_hazard_M~q ),
	.datab(!\M_wr_data_unfiltered[17]~18_combout ),
	.datac(!\E_src2_prelim[17]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_stw_data[17]~35_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_stw_data[17]~35 .extended_lut = "off";
defparam \E_stw_data[17]~35 .lut_mask = 64'h2727272727272727;
defparam \E_stw_data[17]~35 .shared_arith = "off";

cyclonev_lcell_comb \Add8~93 (
	.dataa(!\E_ctrl_alu_subtract~q ),
	.datab(!\E_ctrl_src2_choose_imm~q ),
	.datac(!\E_stw_data[18]~34_combout ),
	.datad(!\E_src2_imm[18]~q ),
	.datae(gnd),
	.dataf(!\E_src1[18]~38_combout ),
	.datag(gnd),
	.cin(\Add8~86 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add8~93_sumout ),
	.cout(\Add8~94 ),
	.shareout());
defparam \Add8~93 .extended_lut = "off";
defparam \Add8~93 .lut_mask = 64'h0000FF0000006996;
defparam \Add8~93 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[18]~32 (
	.dataa(!\E_ctrl_src2_choose_imm~q ),
	.datab(!\E_compare_op[1]~q ),
	.datac(!\E_compare_op[0]~q ),
	.datad(!\E_src1[18]~38_combout ),
	.datae(!\E_src2_imm[18]~q ),
	.dataf(!\E_stw_data[18]~34_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[18]~32_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[18]~32 .extended_lut = "off";
defparam \E_alu_result[18]~32 .lut_mask = 64'h6996966996696996;
defparam \E_alu_result[18]~32 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[18]~33 (
	.dataa(!\E_ctrl_logic~q ),
	.datab(!\E_alu_result~0_combout ),
	.datac(!\Add8~93_sumout ),
	.datad(!\E_alu_result[18]~32_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[18]~33_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[18]~33 .extended_lut = "off";
defparam \E_alu_result[18]~33 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \E_alu_result[18]~33 .shared_arith = "off";

dffeas \M_alu_result[18] (
	.clk(clk_clk),
	.d(\E_alu_result[18]~33_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\M_alu_result[18]~q ),
	.prn(vcc));
defparam \M_alu_result[18] .is_wysiwyg = "true";
defparam \M_alu_result[18] .power_up = "low";

cyclonev_lcell_comb \E_src1[18]~36 (
	.dataa(!\M_ctrl_shift_rot~q ),
	.datab(!\av_ld_or_div_done~q ),
	.datac(!\E_src1_hazard_M~q ),
	.datad(!\M_shift_rot_result[18]~q ),
	.datae(!\av_ld_data_aligned_or_div[18]~q ),
	.dataf(!\M_alu_result[18]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_src1[18]~36_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_src1[18]~36 .extended_lut = "off";
defparam \E_src1[18]~36 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \E_src1[18]~36 .shared_arith = "off";

cyclonev_lcell_comb \D_src1_prelim[18]~20 (
	.dataa(!\M_wr_data_unfiltered[18]~23_combout ),
	.datab(!\D_src1_hazard_M~combout ),
	.datac(!\D_src1_hazard_W~combout ),
	.datad(!\W_wr_data[18]~q ),
	.datae(!\processor_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[18] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_prelim[18]~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src1_prelim[18]~20 .extended_lut = "off";
defparam \D_src1_prelim[18]~20 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \D_src1_prelim[18]~20 .shared_arith = "off";

dffeas \E_src1_prelim[18] (
	.clk(clk_clk),
	.d(\D_src1_prelim[18]~20_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_src1_prelim[18]~q ),
	.prn(vcc));
defparam \E_src1_prelim[18] .is_wysiwyg = "true";
defparam \E_src1_prelim[18] .power_up = "low";

cyclonev_lcell_comb \E_src1[18]~37 (
	.dataa(!\E_src1_hazard_M~q ),
	.datab(!\E_src1_prelim[18]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_src1[18]~37_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_src1[18]~37 .extended_lut = "off";
defparam \E_src1[18]~37 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \E_src1[18]~37 .shared_arith = "off";

cyclonev_lcell_comb \E_src1[18]~38 (
	.dataa(!\E_src1[18]~36_combout ),
	.datab(!\E_src1[18]~37_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_src1[18]~38_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_src1[18]~38 .extended_lut = "off";
defparam \E_src1[18]~38 .lut_mask = 64'h7777777777777777;
defparam \E_src1[18]~38 .shared_arith = "off";

cyclonev_lcell_comb \M_shift_rot_result_nxt[18]~20 (
	.dataa(!\M_shift_rot_stall~q ),
	.datab(!\M_ctrl_shift_rot_right~q ),
	.datac(!\M_shift_rot_result[19]~q ),
	.datad(!\E_src1[18]~38_combout ),
	.datae(!\M_shift_rot_result[17]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_shift_rot_result_nxt[18]~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_shift_rot_result_nxt[18]~20 .extended_lut = "off";
defparam \M_shift_rot_result_nxt[18]~20 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \M_shift_rot_result_nxt[18]~20 .shared_arith = "off";

dffeas \M_shift_rot_result[18] (
	.clk(clk_clk),
	.d(\M_shift_rot_result_nxt[18]~20_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\M_shift_rot_result[18]~q ),
	.prn(vcc));
defparam \M_shift_rot_result[18] .is_wysiwyg = "true";
defparam \M_shift_rot_result[18] .power_up = "low";

dffeas \W_wr_data[19] (
	.clk(clk_clk),
	.d(\M_wr_data_unfiltered[19]~22_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\W_wr_data[19]~q ),
	.prn(vcc));
defparam \W_wr_data[19] .is_wysiwyg = "true";
defparam \W_wr_data[19] .power_up = "low";

cyclonev_lcell_comb \D_src1_prelim[19]~22 (
	.dataa(!\M_wr_data_unfiltered[19]~22_combout ),
	.datab(!\D_src1_hazard_M~combout ),
	.datac(!\D_src1_hazard_W~combout ),
	.datad(!\W_wr_data[19]~q ),
	.datae(!\processor_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[19] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_prelim[19]~22_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src1_prelim[19]~22 .extended_lut = "off";
defparam \D_src1_prelim[19]~22 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \D_src1_prelim[19]~22 .shared_arith = "off";

dffeas \E_src1_prelim[19] (
	.clk(clk_clk),
	.d(\D_src1_prelim[19]~22_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_src1_prelim[19]~q ),
	.prn(vcc));
defparam \E_src1_prelim[19] .is_wysiwyg = "true";
defparam \E_src1_prelim[19] .power_up = "low";

cyclonev_lcell_comb \E_src1[19]~40 (
	.dataa(!\E_src1_hazard_M~q ),
	.datab(!\M_wr_data_unfiltered[19]~22_combout ),
	.datac(!\E_src1_prelim[19]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_src1[19]~40_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_src1[19]~40 .extended_lut = "off";
defparam \E_src1[19]~40 .lut_mask = 64'h2727272727272727;
defparam \E_src1[19]~40 .shared_arith = "off";

cyclonev_lcell_comb \M_shift_rot_result_nxt[19]~22 (
	.dataa(!\M_shift_rot_stall~q ),
	.datab(!\M_ctrl_shift_rot_right~q ),
	.datac(!\M_shift_rot_result[20]~q ),
	.datad(!\M_shift_rot_result[18]~q ),
	.datae(!\E_src1[19]~40_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_shift_rot_result_nxt[19]~22_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_shift_rot_result_nxt[19]~22 .extended_lut = "off";
defparam \M_shift_rot_result_nxt[19]~22 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \M_shift_rot_result_nxt[19]~22 .shared_arith = "off";

dffeas \M_shift_rot_result[19] (
	.clk(clk_clk),
	.d(\M_shift_rot_result_nxt[19]~22_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\M_shift_rot_result[19]~q ),
	.prn(vcc));
defparam \M_shift_rot_result[19] .is_wysiwyg = "true";
defparam \M_shift_rot_result[19] .power_up = "low";

dffeas \av_ld_data_aligned_or_div[19] (
	.clk(clk_clk),
	.d(\av_fill_bit~0_combout ),
	.asdata(\d_readdata_d1[19]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\M_iw[4]~q ),
	.ena(vcc),
	.q(\av_ld_data_aligned_or_div[19]~q ),
	.prn(vcc));
defparam \av_ld_data_aligned_or_div[19] .is_wysiwyg = "true";
defparam \av_ld_data_aligned_or_div[19] .power_up = "low";

dffeas \E_src2_imm[19] (
	.clk(clk_clk),
	.d(\D_iw[21]~q ),
	.asdata(\D_iw[9]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\D_ctrl_unsigned_lo_imm16~combout ),
	.sload(\Equal171~0_combout ),
	.ena(\W_stall~combout ),
	.q(\E_src2_imm[19]~q ),
	.prn(vcc));
defparam \E_src2_imm[19] .is_wysiwyg = "true";
defparam \E_src2_imm[19] .power_up = "low";

cyclonev_lcell_comb \Add8~117 (
	.dataa(!\E_ctrl_alu_subtract~q ),
	.datab(!\E_ctrl_src2_choose_imm~q ),
	.datac(!\E_stw_data[19]~42_combout ),
	.datad(!\E_src2_imm[19]~q ),
	.datae(gnd),
	.dataf(!\E_src1[19]~40_combout ),
	.datag(gnd),
	.cin(\Add8~94 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add8~117_sumout ),
	.cout(\Add8~118 ),
	.shareout());
defparam \Add8~117 .extended_lut = "off";
defparam \Add8~117 .lut_mask = 64'h0000FF0000006996;
defparam \Add8~117 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_prelim[19]~31 (
	.dataa(!\M_wr_data_unfiltered[19]~22_combout ),
	.datab(!\D_src2_hazard_M~combout ),
	.datac(!\D_src2_hazard_W~combout ),
	.datad(!\W_wr_data[19]~q ),
	.datae(!\processor_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[19] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_prelim[19]~31_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_prelim[19]~31 .extended_lut = "off";
defparam \D_src2_prelim[19]~31 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \D_src2_prelim[19]~31 .shared_arith = "off";

dffeas \E_src2_prelim[19] (
	.clk(clk_clk),
	.d(\D_src2_prelim[19]~31_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_src2_prelim[19]~q ),
	.prn(vcc));
defparam \E_src2_prelim[19] .is_wysiwyg = "true";
defparam \E_src2_prelim[19] .power_up = "low";

cyclonev_lcell_comb \E_arith_src2[19]~16 (
	.dataa(!\E_src2_hazard_M~q ),
	.datab(!\E_ctrl_src2_choose_imm~q ),
	.datac(!\M_wr_data_unfiltered[19]~22_combout ),
	.datad(!\E_src2_imm[19]~q ),
	.datae(!\E_src2_prelim[19]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_arith_src2[19]~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_arith_src2[19]~16 .extended_lut = "off";
defparam \E_arith_src2[19]~16 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \E_arith_src2[19]~16 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[19]~46 (
	.dataa(!\E_compare_op[1]~q ),
	.datab(!\E_compare_op[0]~q ),
	.datac(!\E_arith_src2[19]~16_combout ),
	.datad(!\E_src1[19]~40_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[19]~46_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[19]~46 .extended_lut = "off";
defparam \E_alu_result[19]~46 .lut_mask = 64'h6996699669966996;
defparam \E_alu_result[19]~46 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[19]~47 (
	.dataa(!\E_ctrl_logic~q ),
	.datab(!\E_alu_result~0_combout ),
	.datac(!\Add8~117_sumout ),
	.datad(!\E_alu_result[19]~46_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[19]~47_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[19]~47 .extended_lut = "off";
defparam \E_alu_result[19]~47 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \E_alu_result[19]~47 .shared_arith = "off";

dffeas \M_alu_result[19] (
	.clk(clk_clk),
	.d(\E_alu_result[19]~47_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\M_alu_result[19]~q ),
	.prn(vcc));
defparam \M_alu_result[19] .is_wysiwyg = "true";
defparam \M_alu_result[19] .power_up = "low";

cyclonev_lcell_comb \M_wr_data_unfiltered[19]~22 (
	.dataa(!\M_ctrl_shift_rot~q ),
	.datab(!\av_ld_or_div_done~q ),
	.datac(!\M_shift_rot_result[19]~q ),
	.datad(!\av_ld_data_aligned_or_div[19]~q ),
	.datae(!\M_alu_result[19]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_wr_data_unfiltered[19]~22_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_wr_data_unfiltered[19]~22 .extended_lut = "off";
defparam \M_wr_data_unfiltered[19]~22 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \M_wr_data_unfiltered[19]~22 .shared_arith = "off";

cyclonev_lcell_comb \E_stw_data[19]~42 (
	.dataa(!\E_src2_hazard_M~q ),
	.datab(!\M_wr_data_unfiltered[19]~22_combout ),
	.datac(!\E_src2_prelim[19]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_stw_data[19]~42_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_stw_data[19]~42 .extended_lut = "off";
defparam \E_stw_data[19]~42 .lut_mask = 64'h2727272727272727;
defparam \E_stw_data[19]~42 .shared_arith = "off";

cyclonev_lcell_comb \Add8~109 (
	.dataa(!\E_ctrl_alu_subtract~q ),
	.datab(!\E_ctrl_src2_choose_imm~q ),
	.datac(!\E_stw_data[20]~25_combout ),
	.datad(!\E_src2_imm[20]~q ),
	.datae(gnd),
	.dataf(!\E_src1[20]~50_combout ),
	.datag(gnd),
	.cin(\Add8~118 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add8~109_sumout ),
	.cout(\Add8~110 ),
	.shareout());
defparam \Add8~109 .extended_lut = "off";
defparam \Add8~109 .lut_mask = 64'h0000FF0000006996;
defparam \Add8~109 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[20]~40 (
	.dataa(!\E_ctrl_src2_choose_imm~q ),
	.datab(!\E_compare_op[1]~q ),
	.datac(!\E_compare_op[0]~q ),
	.datad(!\E_src1[20]~50_combout ),
	.datae(!\E_src2_imm[20]~q ),
	.dataf(!\E_stw_data[20]~25_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[20]~40_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[20]~40 .extended_lut = "off";
defparam \E_alu_result[20]~40 .lut_mask = 64'h6996966996696996;
defparam \E_alu_result[20]~40 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[20]~41 (
	.dataa(!\E_ctrl_logic~q ),
	.datab(!\E_alu_result~0_combout ),
	.datac(!\Add8~109_sumout ),
	.datad(!\E_alu_result[20]~40_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[20]~41_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[20]~41 .extended_lut = "off";
defparam \E_alu_result[20]~41 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \E_alu_result[20]~41 .shared_arith = "off";

dffeas \M_alu_result[20] (
	.clk(clk_clk),
	.d(\E_alu_result[20]~41_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\M_alu_result[20]~q ),
	.prn(vcc));
defparam \M_alu_result[20] .is_wysiwyg = "true";
defparam \M_alu_result[20] .power_up = "low";

cyclonev_lcell_comb \E_src1[20]~48 (
	.dataa(!\M_ctrl_shift_rot~q ),
	.datab(!\av_ld_or_div_done~q ),
	.datac(!\E_src1_hazard_M~q ),
	.datad(!\M_shift_rot_result[20]~q ),
	.datae(!\av_ld_data_aligned_or_div[20]~q ),
	.dataf(!\M_alu_result[20]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_src1[20]~48_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_src1[20]~48 .extended_lut = "off";
defparam \E_src1[20]~48 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \E_src1[20]~48 .shared_arith = "off";

cyclonev_lcell_comb \D_src1_prelim[20]~26 (
	.dataa(!\M_wr_data_unfiltered[20]~28_combout ),
	.datab(!\D_src1_hazard_M~combout ),
	.datac(!\D_src1_hazard_W~combout ),
	.datad(!\W_wr_data[20]~q ),
	.datae(!\processor_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[20] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_prelim[20]~26_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src1_prelim[20]~26 .extended_lut = "off";
defparam \D_src1_prelim[20]~26 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \D_src1_prelim[20]~26 .shared_arith = "off";

dffeas \E_src1_prelim[20] (
	.clk(clk_clk),
	.d(\D_src1_prelim[20]~26_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_src1_prelim[20]~q ),
	.prn(vcc));
defparam \E_src1_prelim[20] .is_wysiwyg = "true";
defparam \E_src1_prelim[20] .power_up = "low";

cyclonev_lcell_comb \E_src1[20]~49 (
	.dataa(!\E_src1_hazard_M~q ),
	.datab(!\E_src1_prelim[20]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_src1[20]~49_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_src1[20]~49 .extended_lut = "off";
defparam \E_src1[20]~49 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \E_src1[20]~49 .shared_arith = "off";

cyclonev_lcell_comb \E_src1[20]~50 (
	.dataa(!\E_src1[20]~48_combout ),
	.datab(!\E_src1[20]~49_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_src1[20]~50_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_src1[20]~50 .extended_lut = "off";
defparam \E_src1[20]~50 .lut_mask = 64'h7777777777777777;
defparam \E_src1[20]~50 .shared_arith = "off";

cyclonev_lcell_comb \M_shift_rot_result_nxt[20]~26 (
	.dataa(!\M_shift_rot_stall~q ),
	.datab(!\M_ctrl_shift_rot_right~q ),
	.datac(!\M_shift_rot_result[21]~q ),
	.datad(!\E_src1[20]~50_combout ),
	.datae(!\M_shift_rot_result[19]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_shift_rot_result_nxt[20]~26_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_shift_rot_result_nxt[20]~26 .extended_lut = "off";
defparam \M_shift_rot_result_nxt[20]~26 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \M_shift_rot_result_nxt[20]~26 .shared_arith = "off";

dffeas \M_shift_rot_result[20] (
	.clk(clk_clk),
	.d(\M_shift_rot_result_nxt[20]~26_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\M_shift_rot_result[20]~q ),
	.prn(vcc));
defparam \M_shift_rot_result[20] .is_wysiwyg = "true";
defparam \M_shift_rot_result[20] .power_up = "low";

dffeas \W_wr_data[21] (
	.clk(clk_clk),
	.d(\M_wr_data_unfiltered[21]~21_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\W_wr_data[21]~q ),
	.prn(vcc));
defparam \W_wr_data[21] .is_wysiwyg = "true";
defparam \W_wr_data[21] .power_up = "low";

cyclonev_lcell_comb \D_src1_prelim[21]~25 (
	.dataa(!\M_wr_data_unfiltered[21]~21_combout ),
	.datab(!\D_src1_hazard_M~combout ),
	.datac(!\D_src1_hazard_W~combout ),
	.datad(!\W_wr_data[21]~q ),
	.datae(!\processor_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[21] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_prelim[21]~25_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src1_prelim[21]~25 .extended_lut = "off";
defparam \D_src1_prelim[21]~25 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \D_src1_prelim[21]~25 .shared_arith = "off";

dffeas \E_src1_prelim[21] (
	.clk(clk_clk),
	.d(\D_src1_prelim[21]~25_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_src1_prelim[21]~q ),
	.prn(vcc));
defparam \E_src1_prelim[21] .is_wysiwyg = "true";
defparam \E_src1_prelim[21] .power_up = "low";

cyclonev_lcell_comb \E_src1[21]~47 (
	.dataa(!\E_src1_hazard_M~q ),
	.datab(!\M_wr_data_unfiltered[21]~21_combout ),
	.datac(!\E_src1_prelim[21]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_src1[21]~47_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_src1[21]~47 .extended_lut = "off";
defparam \E_src1[21]~47 .lut_mask = 64'h2727272727272727;
defparam \E_src1[21]~47 .shared_arith = "off";

cyclonev_lcell_comb \M_shift_rot_result_nxt[21]~25 (
	.dataa(!\M_shift_rot_stall~q ),
	.datab(!\M_ctrl_shift_rot_right~q ),
	.datac(!\M_shift_rot_result[22]~q ),
	.datad(!\M_shift_rot_result[20]~q ),
	.datae(!\E_src1[21]~47_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_shift_rot_result_nxt[21]~25_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_shift_rot_result_nxt[21]~25 .extended_lut = "off";
defparam \M_shift_rot_result_nxt[21]~25 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \M_shift_rot_result_nxt[21]~25 .shared_arith = "off";

dffeas \M_shift_rot_result[21] (
	.clk(clk_clk),
	.d(\M_shift_rot_result_nxt[21]~25_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\M_shift_rot_result[21]~q ),
	.prn(vcc));
defparam \M_shift_rot_result[21] .is_wysiwyg = "true";
defparam \M_shift_rot_result[21] .power_up = "low";

dffeas \av_ld_data_aligned_or_div[21] (
	.clk(clk_clk),
	.d(\av_fill_bit~0_combout ),
	.asdata(\d_readdata_d1[21]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\M_iw[4]~q ),
	.ena(vcc),
	.q(\av_ld_data_aligned_or_div[21]~q ),
	.prn(vcc));
defparam \av_ld_data_aligned_or_div[21] .is_wysiwyg = "true";
defparam \av_ld_data_aligned_or_div[21] .power_up = "low";

dffeas \E_src2_imm[21] (
	.clk(clk_clk),
	.d(\D_iw[21]~q ),
	.asdata(\D_iw[11]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\D_ctrl_unsigned_lo_imm16~combout ),
	.sload(\Equal171~0_combout ),
	.ena(\W_stall~combout ),
	.q(\E_src2_imm[21]~q ),
	.prn(vcc));
defparam \E_src2_imm[21] .is_wysiwyg = "true";
defparam \E_src2_imm[21] .power_up = "low";

cyclonev_lcell_comb \Add8~105 (
	.dataa(!\E_ctrl_alu_subtract~q ),
	.datab(!\E_ctrl_src2_choose_imm~q ),
	.datac(!\E_stw_data[21]~21_combout ),
	.datad(!\E_src2_imm[21]~q ),
	.datae(gnd),
	.dataf(!\E_src1[21]~47_combout ),
	.datag(gnd),
	.cin(\Add8~110 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add8~105_sumout ),
	.cout(\Add8~106 ),
	.shareout());
defparam \Add8~105 .extended_lut = "off";
defparam \Add8~105 .lut_mask = 64'h0000FF0000006996;
defparam \Add8~105 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_prelim[21]~21 (
	.dataa(!\M_wr_data_unfiltered[21]~21_combout ),
	.datab(!\D_src2_hazard_M~combout ),
	.datac(!\D_src2_hazard_W~combout ),
	.datad(!\W_wr_data[21]~q ),
	.datae(!\processor_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[21] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_prelim[21]~21_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_prelim[21]~21 .extended_lut = "off";
defparam \D_src2_prelim[21]~21 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \D_src2_prelim[21]~21 .shared_arith = "off";

dffeas \E_src2_prelim[21] (
	.clk(clk_clk),
	.d(\D_src2_prelim[21]~21_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_src2_prelim[21]~q ),
	.prn(vcc));
defparam \E_src2_prelim[21] .is_wysiwyg = "true";
defparam \E_src2_prelim[21] .power_up = "low";

cyclonev_lcell_comb \E_arith_src2[21]~15 (
	.dataa(!\E_src2_hazard_M~q ),
	.datab(!\E_ctrl_src2_choose_imm~q ),
	.datac(!\M_wr_data_unfiltered[21]~21_combout ),
	.datad(!\E_src2_imm[21]~q ),
	.datae(!\E_src2_prelim[21]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_arith_src2[21]~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_arith_src2[21]~15 .extended_lut = "off";
defparam \E_arith_src2[21]~15 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \E_arith_src2[21]~15 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[21]~38 (
	.dataa(!\E_compare_op[1]~q ),
	.datab(!\E_compare_op[0]~q ),
	.datac(!\E_arith_src2[21]~15_combout ),
	.datad(!\E_src1[21]~47_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[21]~38_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[21]~38 .extended_lut = "off";
defparam \E_alu_result[21]~38 .lut_mask = 64'h6996699669966996;
defparam \E_alu_result[21]~38 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[21]~39 (
	.dataa(!\E_ctrl_logic~q ),
	.datab(!\E_alu_result~0_combout ),
	.datac(!\Add8~105_sumout ),
	.datad(!\E_alu_result[21]~38_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[21]~39_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[21]~39 .extended_lut = "off";
defparam \E_alu_result[21]~39 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \E_alu_result[21]~39 .shared_arith = "off";

dffeas \M_alu_result[21] (
	.clk(clk_clk),
	.d(\E_alu_result[21]~39_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\M_alu_result[21]~q ),
	.prn(vcc));
defparam \M_alu_result[21] .is_wysiwyg = "true";
defparam \M_alu_result[21] .power_up = "low";

cyclonev_lcell_comb \M_wr_data_unfiltered[21]~21 (
	.dataa(!\M_ctrl_shift_rot~q ),
	.datab(!\av_ld_or_div_done~q ),
	.datac(!\M_shift_rot_result[21]~q ),
	.datad(!\av_ld_data_aligned_or_div[21]~q ),
	.datae(!\M_alu_result[21]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_wr_data_unfiltered[21]~21_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_wr_data_unfiltered[21]~21 .extended_lut = "off";
defparam \M_wr_data_unfiltered[21]~21 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \M_wr_data_unfiltered[21]~21 .shared_arith = "off";

cyclonev_lcell_comb \E_stw_data[21]~21 (
	.dataa(!\E_src2_hazard_M~q ),
	.datab(!\M_wr_data_unfiltered[21]~21_combout ),
	.datac(!\E_src2_prelim[21]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_stw_data[21]~21_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_stw_data[21]~21 .extended_lut = "off";
defparam \E_stw_data[21]~21 .lut_mask = 64'h2727272727272727;
defparam \E_stw_data[21]~21 .shared_arith = "off";

cyclonev_lcell_comb \Add8~113 (
	.dataa(!\E_ctrl_alu_subtract~q ),
	.datab(!\E_ctrl_src2_choose_imm~q ),
	.datac(!\E_stw_data[22]~31_combout ),
	.datad(!\E_src2_imm[22]~q ),
	.datae(gnd),
	.dataf(!\E_src1[22]~53_combout ),
	.datag(gnd),
	.cin(\Add8~106 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add8~113_sumout ),
	.cout(\Add8~114 ),
	.shareout());
defparam \Add8~113 .extended_lut = "off";
defparam \Add8~113 .lut_mask = 64'h0000FF0000006996;
defparam \Add8~113 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[22]~44 (
	.dataa(!\E_ctrl_src2_choose_imm~q ),
	.datab(!\E_compare_op[1]~q ),
	.datac(!\E_compare_op[0]~q ),
	.datad(!\E_src1[22]~53_combout ),
	.datae(!\E_src2_imm[22]~q ),
	.dataf(!\E_stw_data[22]~31_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[22]~44_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[22]~44 .extended_lut = "off";
defparam \E_alu_result[22]~44 .lut_mask = 64'h6996966996696996;
defparam \E_alu_result[22]~44 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[22]~45 (
	.dataa(!\E_ctrl_logic~q ),
	.datab(!\E_alu_result~0_combout ),
	.datac(!\Add8~113_sumout ),
	.datad(!\E_alu_result[22]~44_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[22]~45_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[22]~45 .extended_lut = "off";
defparam \E_alu_result[22]~45 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \E_alu_result[22]~45 .shared_arith = "off";

dffeas \M_alu_result[22] (
	.clk(clk_clk),
	.d(\E_alu_result[22]~45_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\M_alu_result[22]~q ),
	.prn(vcc));
defparam \M_alu_result[22] .is_wysiwyg = "true";
defparam \M_alu_result[22] .power_up = "low";

cyclonev_lcell_comb \E_src1[22]~51 (
	.dataa(!\M_ctrl_shift_rot~q ),
	.datab(!\av_ld_or_div_done~q ),
	.datac(!\E_src1_hazard_M~q ),
	.datad(!\M_shift_rot_result[22]~q ),
	.datae(!\av_ld_data_aligned_or_div[22]~q ),
	.dataf(!\M_alu_result[22]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_src1[22]~51_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_src1[22]~51 .extended_lut = "off";
defparam \E_src1[22]~51 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \E_src1[22]~51 .shared_arith = "off";

cyclonev_lcell_comb \D_src1_prelim[22]~27 (
	.dataa(!\M_wr_data_unfiltered[22]~30_combout ),
	.datab(!\D_src1_hazard_M~combout ),
	.datac(!\D_src1_hazard_W~combout ),
	.datad(!\W_wr_data[22]~q ),
	.datae(!\processor_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[22] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_prelim[22]~27_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src1_prelim[22]~27 .extended_lut = "off";
defparam \D_src1_prelim[22]~27 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \D_src1_prelim[22]~27 .shared_arith = "off";

dffeas \E_src1_prelim[22] (
	.clk(clk_clk),
	.d(\D_src1_prelim[22]~27_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_src1_prelim[22]~q ),
	.prn(vcc));
defparam \E_src1_prelim[22] .is_wysiwyg = "true";
defparam \E_src1_prelim[22] .power_up = "low";

cyclonev_lcell_comb \E_src1[22]~52 (
	.dataa(!\E_src1_hazard_M~q ),
	.datab(!\E_src1_prelim[22]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_src1[22]~52_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_src1[22]~52 .extended_lut = "off";
defparam \E_src1[22]~52 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \E_src1[22]~52 .shared_arith = "off";

cyclonev_lcell_comb \E_src1[22]~53 (
	.dataa(!\E_src1[22]~51_combout ),
	.datab(!\E_src1[22]~52_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_src1[22]~53_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_src1[22]~53 .extended_lut = "off";
defparam \E_src1[22]~53 .lut_mask = 64'h7777777777777777;
defparam \E_src1[22]~53 .shared_arith = "off";

cyclonev_lcell_comb \M_shift_rot_result_nxt[22]~27 (
	.dataa(!\M_shift_rot_stall~q ),
	.datab(!\M_ctrl_shift_rot_right~q ),
	.datac(!\M_shift_rot_result[23]~q ),
	.datad(!\E_src1[22]~53_combout ),
	.datae(!\M_shift_rot_result[21]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_shift_rot_result_nxt[22]~27_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_shift_rot_result_nxt[22]~27 .extended_lut = "off";
defparam \M_shift_rot_result_nxt[22]~27 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \M_shift_rot_result_nxt[22]~27 .shared_arith = "off";

dffeas \M_shift_rot_result[22] (
	.clk(clk_clk),
	.d(\M_shift_rot_result_nxt[22]~27_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\M_shift_rot_result[22]~q ),
	.prn(vcc));
defparam \M_shift_rot_result[22] .is_wysiwyg = "true";
defparam \M_shift_rot_result[22] .power_up = "low";

dffeas \W_wr_data[23] (
	.clk(clk_clk),
	.d(\M_wr_data_unfiltered[23]~24_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\W_wr_data[23]~q ),
	.prn(vcc));
defparam \W_wr_data[23] .is_wysiwyg = "true";
defparam \W_wr_data[23] .power_up = "low";

cyclonev_lcell_comb \D_src1_prelim[23]~28 (
	.dataa(!\M_wr_data_unfiltered[23]~24_combout ),
	.datab(!\D_src1_hazard_M~combout ),
	.datac(!\D_src1_hazard_W~combout ),
	.datad(!\W_wr_data[23]~q ),
	.datae(!\processor_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[23] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_prelim[23]~28_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src1_prelim[23]~28 .extended_lut = "off";
defparam \D_src1_prelim[23]~28 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \D_src1_prelim[23]~28 .shared_arith = "off";

dffeas \E_src1_prelim[23] (
	.clk(clk_clk),
	.d(\D_src1_prelim[23]~28_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_src1_prelim[23]~q ),
	.prn(vcc));
defparam \E_src1_prelim[23] .is_wysiwyg = "true";
defparam \E_src1_prelim[23] .power_up = "low";

cyclonev_lcell_comb \E_src1[23]~54 (
	.dataa(!\E_src1_hazard_M~q ),
	.datab(!\M_wr_data_unfiltered[23]~24_combout ),
	.datac(!\E_src1_prelim[23]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_src1[23]~54_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_src1[23]~54 .extended_lut = "off";
defparam \E_src1[23]~54 .lut_mask = 64'h2727272727272727;
defparam \E_src1[23]~54 .shared_arith = "off";

cyclonev_lcell_comb \M_shift_rot_result_nxt[23]~28 (
	.dataa(!\M_shift_rot_stall~q ),
	.datab(!\M_ctrl_shift_rot_right~q ),
	.datac(!\M_shift_rot_result[24]~q ),
	.datad(!\M_shift_rot_result[22]~q ),
	.datae(!\E_src1[23]~54_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_shift_rot_result_nxt[23]~28_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_shift_rot_result_nxt[23]~28 .extended_lut = "off";
defparam \M_shift_rot_result_nxt[23]~28 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \M_shift_rot_result_nxt[23]~28 .shared_arith = "off";

dffeas \M_shift_rot_result[23] (
	.clk(clk_clk),
	.d(\M_shift_rot_result_nxt[23]~28_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\M_shift_rot_result[23]~q ),
	.prn(vcc));
defparam \M_shift_rot_result[23] .is_wysiwyg = "true";
defparam \M_shift_rot_result[23] .power_up = "low";

dffeas \av_ld_data_aligned_or_div[23] (
	.clk(clk_clk),
	.d(\av_fill_bit~0_combout ),
	.asdata(\d_readdata_d1[23]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\M_iw[4]~q ),
	.ena(vcc),
	.q(\av_ld_data_aligned_or_div[23]~q ),
	.prn(vcc));
defparam \av_ld_data_aligned_or_div[23] .is_wysiwyg = "true";
defparam \av_ld_data_aligned_or_div[23] .power_up = "low";

dffeas \E_src2_imm[23] (
	.clk(clk_clk),
	.d(\D_iw[21]~q ),
	.asdata(\D_iw[13]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\D_ctrl_unsigned_lo_imm16~combout ),
	.sload(\Equal171~0_combout ),
	.ena(\W_stall~combout ),
	.q(\E_src2_imm[23]~q ),
	.prn(vcc));
defparam \E_src2_imm[23] .is_wysiwyg = "true";
defparam \E_src2_imm[23] .power_up = "low";

cyclonev_lcell_comb \Add8~121 (
	.dataa(!\E_ctrl_alu_subtract~q ),
	.datab(!\E_ctrl_src2_choose_imm~q ),
	.datac(!\E_stw_data[23]~36_combout ),
	.datad(!\E_src2_imm[23]~q ),
	.datae(gnd),
	.dataf(!\E_src1[23]~54_combout ),
	.datag(gnd),
	.cin(\Add8~114 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add8~121_sumout ),
	.cout(\Add8~122 ),
	.shareout());
defparam \Add8~121 .extended_lut = "off";
defparam \Add8~121 .lut_mask = 64'h0000FF0000006996;
defparam \Add8~121 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_prelim[23]~27 (
	.dataa(!\M_wr_data_unfiltered[23]~24_combout ),
	.datab(!\D_src2_hazard_M~combout ),
	.datac(!\D_src2_hazard_W~combout ),
	.datad(!\W_wr_data[23]~q ),
	.datae(!\processor_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[23] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_prelim[23]~27_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_prelim[23]~27 .extended_lut = "off";
defparam \D_src2_prelim[23]~27 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \D_src2_prelim[23]~27 .shared_arith = "off";

dffeas \E_src2_prelim[23] (
	.clk(clk_clk),
	.d(\D_src2_prelim[23]~27_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_src2_prelim[23]~q ),
	.prn(vcc));
defparam \E_src2_prelim[23] .is_wysiwyg = "true";
defparam \E_src2_prelim[23] .power_up = "low";

cyclonev_lcell_comb \E_arith_src2[23]~17 (
	.dataa(!\E_src2_hazard_M~q ),
	.datab(!\E_ctrl_src2_choose_imm~q ),
	.datac(!\M_wr_data_unfiltered[23]~24_combout ),
	.datad(!\E_src2_imm[23]~q ),
	.datae(!\E_src2_prelim[23]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_arith_src2[23]~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_arith_src2[23]~17 .extended_lut = "off";
defparam \E_arith_src2[23]~17 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \E_arith_src2[23]~17 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[23]~48 (
	.dataa(!\E_compare_op[1]~q ),
	.datab(!\E_compare_op[0]~q ),
	.datac(!\E_arith_src2[23]~17_combout ),
	.datad(!\E_src1[23]~54_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[23]~48_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[23]~48 .extended_lut = "off";
defparam \E_alu_result[23]~48 .lut_mask = 64'h6996699669966996;
defparam \E_alu_result[23]~48 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[23]~49 (
	.dataa(!\E_ctrl_logic~q ),
	.datab(!\E_alu_result~0_combout ),
	.datac(!\Add8~121_sumout ),
	.datad(!\E_alu_result[23]~48_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[23]~49_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[23]~49 .extended_lut = "off";
defparam \E_alu_result[23]~49 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \E_alu_result[23]~49 .shared_arith = "off";

dffeas \M_alu_result[23] (
	.clk(clk_clk),
	.d(\E_alu_result[23]~49_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\M_alu_result[23]~q ),
	.prn(vcc));
defparam \M_alu_result[23] .is_wysiwyg = "true";
defparam \M_alu_result[23] .power_up = "low";

cyclonev_lcell_comb \M_wr_data_unfiltered[23]~24 (
	.dataa(!\M_ctrl_shift_rot~q ),
	.datab(!\av_ld_or_div_done~q ),
	.datac(!\M_shift_rot_result[23]~q ),
	.datad(!\av_ld_data_aligned_or_div[23]~q ),
	.datae(!\M_alu_result[23]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_wr_data_unfiltered[23]~24_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_wr_data_unfiltered[23]~24 .extended_lut = "off";
defparam \M_wr_data_unfiltered[23]~24 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \M_wr_data_unfiltered[23]~24 .shared_arith = "off";

cyclonev_lcell_comb \E_stw_data[23]~36 (
	.dataa(!\E_src2_hazard_M~q ),
	.datab(!\M_wr_data_unfiltered[23]~24_combout ),
	.datac(!\E_src2_prelim[23]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_stw_data[23]~36_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_stw_data[23]~36 .extended_lut = "off";
defparam \E_stw_data[23]~36 .lut_mask = 64'h2727272727272727;
defparam \E_stw_data[23]~36 .shared_arith = "off";

cyclonev_lcell_comb \Add8~97 (
	.dataa(!\E_ctrl_alu_subtract~q ),
	.datab(!\E_ctrl_src2_choose_imm~q ),
	.datac(!\E_stw_data[24]~20_combout ),
	.datad(!\E_src2_imm[24]~q ),
	.datae(gnd),
	.dataf(!\E_src1[24]~46_combout ),
	.datag(gnd),
	.cin(\Add8~122 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add8~97_sumout ),
	.cout(\Add8~98 ),
	.shareout());
defparam \Add8~97 .extended_lut = "off";
defparam \Add8~97 .lut_mask = 64'h0000FF0000006996;
defparam \Add8~97 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[24]~36 (
	.dataa(!\E_ctrl_src2_choose_imm~q ),
	.datab(!\E_compare_op[1]~q ),
	.datac(!\E_compare_op[0]~q ),
	.datad(!\E_src1[24]~46_combout ),
	.datae(!\E_src2_imm[24]~q ),
	.dataf(!\E_stw_data[24]~20_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[24]~36_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[24]~36 .extended_lut = "off";
defparam \E_alu_result[24]~36 .lut_mask = 64'h6996966996696996;
defparam \E_alu_result[24]~36 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[24]~37 (
	.dataa(!\E_ctrl_logic~q ),
	.datab(!\E_alu_result~0_combout ),
	.datac(!\Add8~97_sumout ),
	.datad(!\E_alu_result[24]~36_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[24]~37_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[24]~37 .extended_lut = "off";
defparam \E_alu_result[24]~37 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \E_alu_result[24]~37 .shared_arith = "off";

dffeas \M_alu_result[24] (
	.clk(clk_clk),
	.d(\E_alu_result[24]~37_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\M_alu_result[24]~q ),
	.prn(vcc));
defparam \M_alu_result[24] .is_wysiwyg = "true";
defparam \M_alu_result[24] .power_up = "low";

cyclonev_lcell_comb \E_src1[24]~44 (
	.dataa(!\M_ctrl_shift_rot~q ),
	.datab(!\av_ld_or_div_done~q ),
	.datac(!\E_src1_hazard_M~q ),
	.datad(!\M_shift_rot_result[24]~q ),
	.datae(!\av_ld_data_aligned_or_div[24]~q ),
	.dataf(!\M_alu_result[24]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_src1[24]~44_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_src1[24]~44 .extended_lut = "off";
defparam \E_src1[24]~44 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \E_src1[24]~44 .shared_arith = "off";

cyclonev_lcell_comb \D_src1_prelim[24]~24 (
	.dataa(!\M_wr_data_unfiltered[24]~27_combout ),
	.datab(!\D_src1_hazard_M~combout ),
	.datac(!\D_src1_hazard_W~combout ),
	.datad(!\W_wr_data[24]~q ),
	.datae(!\processor_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[24] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_prelim[24]~24_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src1_prelim[24]~24 .extended_lut = "off";
defparam \D_src1_prelim[24]~24 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \D_src1_prelim[24]~24 .shared_arith = "off";

dffeas \E_src1_prelim[24] (
	.clk(clk_clk),
	.d(\D_src1_prelim[24]~24_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_src1_prelim[24]~q ),
	.prn(vcc));
defparam \E_src1_prelim[24] .is_wysiwyg = "true";
defparam \E_src1_prelim[24] .power_up = "low";

cyclonev_lcell_comb \E_src1[24]~45 (
	.dataa(!\E_src1_hazard_M~q ),
	.datab(!\E_src1_prelim[24]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_src1[24]~45_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_src1[24]~45 .extended_lut = "off";
defparam \E_src1[24]~45 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \E_src1[24]~45 .shared_arith = "off";

cyclonev_lcell_comb \E_src1[24]~46 (
	.dataa(!\E_src1[24]~44_combout ),
	.datab(!\E_src1[24]~45_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_src1[24]~46_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_src1[24]~46 .extended_lut = "off";
defparam \E_src1[24]~46 .lut_mask = 64'h7777777777777777;
defparam \E_src1[24]~46 .shared_arith = "off";

cyclonev_lcell_comb \M_shift_rot_result_nxt[24]~24 (
	.dataa(!\M_shift_rot_stall~q ),
	.datab(!\M_ctrl_shift_rot_right~q ),
	.datac(!\M_shift_rot_result[25]~q ),
	.datad(!\E_src1[24]~46_combout ),
	.datae(!\M_shift_rot_result[23]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_shift_rot_result_nxt[24]~24_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_shift_rot_result_nxt[24]~24 .extended_lut = "off";
defparam \M_shift_rot_result_nxt[24]~24 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \M_shift_rot_result_nxt[24]~24 .shared_arith = "off";

dffeas \M_shift_rot_result[24] (
	.clk(clk_clk),
	.d(\M_shift_rot_result_nxt[24]~24_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\M_shift_rot_result[24]~q ),
	.prn(vcc));
defparam \M_shift_rot_result[24] .is_wysiwyg = "true";
defparam \M_shift_rot_result[24] .power_up = "low";

dffeas \W_wr_data[25] (
	.clk(clk_clk),
	.d(\M_wr_data_unfiltered[25]~26_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\W_wr_data[25]~q ),
	.prn(vcc));
defparam \W_wr_data[25] .is_wysiwyg = "true";
defparam \W_wr_data[25] .power_up = "low";

cyclonev_lcell_comb \D_src1_prelim[25]~31 (
	.dataa(!\M_wr_data_unfiltered[25]~26_combout ),
	.datab(!\D_src1_hazard_M~combout ),
	.datac(!\D_src1_hazard_W~combout ),
	.datad(!\W_wr_data[25]~q ),
	.datae(!\processor_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[25] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_prelim[25]~31_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src1_prelim[25]~31 .extended_lut = "off";
defparam \D_src1_prelim[25]~31 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \D_src1_prelim[25]~31 .shared_arith = "off";

dffeas \E_src1_prelim[25] (
	.clk(clk_clk),
	.d(\D_src1_prelim[25]~31_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_src1_prelim[25]~q ),
	.prn(vcc));
defparam \E_src1_prelim[25] .is_wysiwyg = "true";
defparam \E_src1_prelim[25] .power_up = "low";

cyclonev_lcell_comb \E_src1[25]~59 (
	.dataa(!\E_src1_hazard_M~q ),
	.datab(!\M_wr_data_unfiltered[25]~26_combout ),
	.datac(!\E_src1_prelim[25]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_src1[25]~59_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_src1[25]~59 .extended_lut = "off";
defparam \E_src1[25]~59 .lut_mask = 64'h2727272727272727;
defparam \E_src1[25]~59 .shared_arith = "off";

cyclonev_lcell_comb \M_shift_rot_result_nxt[25]~31 (
	.dataa(!\M_shift_rot_stall~q ),
	.datab(!\M_ctrl_shift_rot_right~q ),
	.datac(!\M_shift_rot_result[26]~q ),
	.datad(!\M_shift_rot_result[24]~q ),
	.datae(!\E_src1[25]~59_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_shift_rot_result_nxt[25]~31_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_shift_rot_result_nxt[25]~31 .extended_lut = "off";
defparam \M_shift_rot_result_nxt[25]~31 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \M_shift_rot_result_nxt[25]~31 .shared_arith = "off";

dffeas \M_shift_rot_result[25] (
	.clk(clk_clk),
	.d(\M_shift_rot_result_nxt[25]~31_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\M_shift_rot_result[25]~q ),
	.prn(vcc));
defparam \M_shift_rot_result[25] .is_wysiwyg = "true";
defparam \M_shift_rot_result[25] .power_up = "low";

dffeas \av_ld_data_aligned_or_div[25] (
	.clk(clk_clk),
	.d(\av_fill_bit~0_combout ),
	.asdata(\d_readdata_d1[25]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\M_iw[4]~q ),
	.ena(vcc),
	.q(\av_ld_data_aligned_or_div[25]~q ),
	.prn(vcc));
defparam \av_ld_data_aligned_or_div[25] .is_wysiwyg = "true";
defparam \av_ld_data_aligned_or_div[25] .power_up = "low";

dffeas \E_src2_imm[25] (
	.clk(clk_clk),
	.d(\D_iw[21]~q ),
	.asdata(\D_iw[15]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\D_ctrl_unsigned_lo_imm16~combout ),
	.sload(\Equal171~0_combout ),
	.ena(\W_stall~combout ),
	.q(\E_src2_imm[25]~q ),
	.prn(vcc));
defparam \E_src2_imm[25] .is_wysiwyg = "true";
defparam \E_src2_imm[25] .power_up = "low";

cyclonev_lcell_comb \Add8~133 (
	.dataa(!\E_ctrl_alu_subtract~q ),
	.datab(!\E_ctrl_src2_choose_imm~q ),
	.datac(!\E_stw_data[25]~41_combout ),
	.datad(!\E_src2_imm[25]~q ),
	.datae(gnd),
	.dataf(!\E_src1[25]~59_combout ),
	.datag(gnd),
	.cin(\Add8~98 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add8~133_sumout ),
	.cout(\Add8~134 ),
	.shareout());
defparam \Add8~133 .extended_lut = "off";
defparam \Add8~133 .lut_mask = 64'h0000FF0000006996;
defparam \Add8~133 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_prelim[25]~30 (
	.dataa(!\M_wr_data_unfiltered[25]~26_combout ),
	.datab(!\D_src2_hazard_M~combout ),
	.datac(!\D_src2_hazard_W~combout ),
	.datad(!\W_wr_data[25]~q ),
	.datae(!\processor_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[25] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_prelim[25]~30_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_prelim[25]~30 .extended_lut = "off";
defparam \D_src2_prelim[25]~30 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \D_src2_prelim[25]~30 .shared_arith = "off";

dffeas \E_src2_prelim[25] (
	.clk(clk_clk),
	.d(\D_src2_prelim[25]~30_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_src2_prelim[25]~q ),
	.prn(vcc));
defparam \E_src2_prelim[25] .is_wysiwyg = "true";
defparam \E_src2_prelim[25] .power_up = "low";

cyclonev_lcell_comb \E_arith_src2[25]~19 (
	.dataa(!\E_src2_hazard_M~q ),
	.datab(!\E_ctrl_src2_choose_imm~q ),
	.datac(!\M_wr_data_unfiltered[25]~26_combout ),
	.datad(!\E_src2_imm[25]~q ),
	.datae(!\E_src2_prelim[25]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_arith_src2[25]~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_arith_src2[25]~19 .extended_lut = "off";
defparam \E_arith_src2[25]~19 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \E_arith_src2[25]~19 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[25]~54 (
	.dataa(!\E_compare_op[1]~q ),
	.datab(!\E_compare_op[0]~q ),
	.datac(!\E_arith_src2[25]~19_combout ),
	.datad(!\E_src1[25]~59_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[25]~54_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[25]~54 .extended_lut = "off";
defparam \E_alu_result[25]~54 .lut_mask = 64'h6996699669966996;
defparam \E_alu_result[25]~54 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[25]~55 (
	.dataa(!\E_ctrl_logic~q ),
	.datab(!\E_alu_result~0_combout ),
	.datac(!\Add8~133_sumout ),
	.datad(!\E_alu_result[25]~54_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[25]~55_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[25]~55 .extended_lut = "off";
defparam \E_alu_result[25]~55 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \E_alu_result[25]~55 .shared_arith = "off";

dffeas \M_alu_result[25] (
	.clk(clk_clk),
	.d(\E_alu_result[25]~55_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\M_alu_result[25]~q ),
	.prn(vcc));
defparam \M_alu_result[25] .is_wysiwyg = "true";
defparam \M_alu_result[25] .power_up = "low";

cyclonev_lcell_comb \M_wr_data_unfiltered[25]~26 (
	.dataa(!\M_ctrl_shift_rot~q ),
	.datab(!\av_ld_or_div_done~q ),
	.datac(!\M_shift_rot_result[25]~q ),
	.datad(!\av_ld_data_aligned_or_div[25]~q ),
	.datae(!\M_alu_result[25]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_wr_data_unfiltered[25]~26_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_wr_data_unfiltered[25]~26 .extended_lut = "off";
defparam \M_wr_data_unfiltered[25]~26 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \M_wr_data_unfiltered[25]~26 .shared_arith = "off";

cyclonev_lcell_comb \E_stw_data[25]~41 (
	.dataa(!\E_src2_hazard_M~q ),
	.datab(!\M_wr_data_unfiltered[25]~26_combout ),
	.datac(!\E_src2_prelim[25]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_stw_data[25]~41_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_stw_data[25]~41 .extended_lut = "off";
defparam \E_stw_data[25]~41 .lut_mask = 64'h2727272727272727;
defparam \E_stw_data[25]~41 .shared_arith = "off";

cyclonev_lcell_comb \Add8~129 (
	.dataa(!\E_ctrl_alu_subtract~q ),
	.datab(!\E_ctrl_src2_choose_imm~q ),
	.datac(!\E_stw_data[26]~40_combout ),
	.datad(!\E_src2_imm[26]~q ),
	.datae(gnd),
	.dataf(!\E_src1[26]~58_combout ),
	.datag(gnd),
	.cin(\Add8~134 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add8~129_sumout ),
	.cout(\Add8~130 ),
	.shareout());
defparam \Add8~129 .extended_lut = "off";
defparam \Add8~129 .lut_mask = 64'h0000FF0000006996;
defparam \Add8~129 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[26]~52 (
	.dataa(!\E_ctrl_src2_choose_imm~q ),
	.datab(!\E_compare_op[1]~q ),
	.datac(!\E_compare_op[0]~q ),
	.datad(!\E_src1[26]~58_combout ),
	.datae(!\E_src2_imm[26]~q ),
	.dataf(!\E_stw_data[26]~40_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[26]~52_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[26]~52 .extended_lut = "off";
defparam \E_alu_result[26]~52 .lut_mask = 64'h6996966996696996;
defparam \E_alu_result[26]~52 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[26]~53 (
	.dataa(!\E_ctrl_logic~q ),
	.datab(!\E_alu_result~0_combout ),
	.datac(!\Add8~129_sumout ),
	.datad(!\E_alu_result[26]~52_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[26]~53_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[26]~53 .extended_lut = "off";
defparam \E_alu_result[26]~53 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \E_alu_result[26]~53 .shared_arith = "off";

dffeas \M_alu_result[26] (
	.clk(clk_clk),
	.d(\E_alu_result[26]~53_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\M_alu_result[26]~q ),
	.prn(vcc));
defparam \M_alu_result[26] .is_wysiwyg = "true";
defparam \M_alu_result[26] .power_up = "low";

cyclonev_lcell_comb \E_src1[26]~56 (
	.dataa(!\M_ctrl_shift_rot~q ),
	.datab(!\av_ld_or_div_done~q ),
	.datac(!\E_src1_hazard_M~q ),
	.datad(!\M_shift_rot_result[26]~q ),
	.datae(!\av_ld_data_aligned_or_div[26]~q ),
	.dataf(!\M_alu_result[26]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_src1[26]~56_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_src1[26]~56 .extended_lut = "off";
defparam \E_src1[26]~56 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \E_src1[26]~56 .shared_arith = "off";

cyclonev_lcell_comb \D_src1_prelim[26]~30 (
	.dataa(!\M_wr_data_unfiltered[26]~31_combout ),
	.datab(!\D_src1_hazard_M~combout ),
	.datac(!\D_src1_hazard_W~combout ),
	.datad(!\W_wr_data[26]~q ),
	.datae(!\processor_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[26] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_prelim[26]~30_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src1_prelim[26]~30 .extended_lut = "off";
defparam \D_src1_prelim[26]~30 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \D_src1_prelim[26]~30 .shared_arith = "off";

dffeas \E_src1_prelim[26] (
	.clk(clk_clk),
	.d(\D_src1_prelim[26]~30_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_src1_prelim[26]~q ),
	.prn(vcc));
defparam \E_src1_prelim[26] .is_wysiwyg = "true";
defparam \E_src1_prelim[26] .power_up = "low";

cyclonev_lcell_comb \E_src1[26]~57 (
	.dataa(!\E_src1_hazard_M~q ),
	.datab(!\E_src1_prelim[26]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_src1[26]~57_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_src1[26]~57 .extended_lut = "off";
defparam \E_src1[26]~57 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \E_src1[26]~57 .shared_arith = "off";

cyclonev_lcell_comb \E_src1[26]~58 (
	.dataa(!\E_src1[26]~56_combout ),
	.datab(!\E_src1[26]~57_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_src1[26]~58_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_src1[26]~58 .extended_lut = "off";
defparam \E_src1[26]~58 .lut_mask = 64'h7777777777777777;
defparam \E_src1[26]~58 .shared_arith = "off";

cyclonev_lcell_comb \M_shift_rot_result_nxt[26]~30 (
	.dataa(!\M_shift_rot_stall~q ),
	.datab(!\M_ctrl_shift_rot_right~q ),
	.datac(!\M_shift_rot_result[27]~q ),
	.datad(!\E_src1[26]~58_combout ),
	.datae(!\M_shift_rot_result[25]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_shift_rot_result_nxt[26]~30_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_shift_rot_result_nxt[26]~30 .extended_lut = "off";
defparam \M_shift_rot_result_nxt[26]~30 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \M_shift_rot_result_nxt[26]~30 .shared_arith = "off";

dffeas \M_shift_rot_result[26] (
	.clk(clk_clk),
	.d(\M_shift_rot_result_nxt[26]~30_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\M_shift_rot_result[26]~q ),
	.prn(vcc));
defparam \M_shift_rot_result[26] .is_wysiwyg = "true";
defparam \M_shift_rot_result[26] .power_up = "low";

dffeas \W_wr_data[27] (
	.clk(clk_clk),
	.d(\M_wr_data_unfiltered[27]~25_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\W_wr_data[27]~q ),
	.prn(vcc));
defparam \W_wr_data[27] .is_wysiwyg = "true";
defparam \W_wr_data[27] .power_up = "low";

cyclonev_lcell_comb \D_src1_prelim[27]~29 (
	.dataa(!\M_wr_data_unfiltered[27]~25_combout ),
	.datab(!\D_src1_hazard_M~combout ),
	.datac(!\D_src1_hazard_W~combout ),
	.datad(!\W_wr_data[27]~q ),
	.datae(!\processor_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[27] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_prelim[27]~29_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src1_prelim[27]~29 .extended_lut = "off";
defparam \D_src1_prelim[27]~29 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \D_src1_prelim[27]~29 .shared_arith = "off";

dffeas \E_src1_prelim[27] (
	.clk(clk_clk),
	.d(\D_src1_prelim[27]~29_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_src1_prelim[27]~q ),
	.prn(vcc));
defparam \E_src1_prelim[27] .is_wysiwyg = "true";
defparam \E_src1_prelim[27] .power_up = "low";

cyclonev_lcell_comb \E_src1[27]~55 (
	.dataa(!\E_src1_hazard_M~q ),
	.datab(!\M_wr_data_unfiltered[27]~25_combout ),
	.datac(!\E_src1_prelim[27]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_src1[27]~55_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_src1[27]~55 .extended_lut = "off";
defparam \E_src1[27]~55 .lut_mask = 64'h2727272727272727;
defparam \E_src1[27]~55 .shared_arith = "off";

cyclonev_lcell_comb \M_shift_rot_result_nxt[27]~29 (
	.dataa(!\M_shift_rot_stall~q ),
	.datab(!\M_ctrl_shift_rot_right~q ),
	.datac(!\M_shift_rot_result[28]~q ),
	.datad(!\M_shift_rot_result[26]~q ),
	.datae(!\E_src1[27]~55_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_shift_rot_result_nxt[27]~29_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_shift_rot_result_nxt[27]~29 .extended_lut = "off";
defparam \M_shift_rot_result_nxt[27]~29 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \M_shift_rot_result_nxt[27]~29 .shared_arith = "off";

dffeas \M_shift_rot_result[27] (
	.clk(clk_clk),
	.d(\M_shift_rot_result_nxt[27]~29_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\M_shift_rot_result[27]~q ),
	.prn(vcc));
defparam \M_shift_rot_result[27] .is_wysiwyg = "true";
defparam \M_shift_rot_result[27] .power_up = "low";

dffeas \av_ld_data_aligned_or_div[27] (
	.clk(clk_clk),
	.d(\av_fill_bit~0_combout ),
	.asdata(\d_readdata_d1[27]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\M_iw[4]~q ),
	.ena(vcc),
	.q(\av_ld_data_aligned_or_div[27]~q ),
	.prn(vcc));
defparam \av_ld_data_aligned_or_div[27] .is_wysiwyg = "true";
defparam \av_ld_data_aligned_or_div[27] .power_up = "low";

dffeas \E_src2_imm[27] (
	.clk(clk_clk),
	.d(\D_iw[21]~q ),
	.asdata(\D_iw[17]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\D_ctrl_unsigned_lo_imm16~combout ),
	.sload(\Equal171~0_combout ),
	.ena(\W_stall~combout ),
	.q(\E_src2_imm[27]~q ),
	.prn(vcc));
defparam \E_src2_imm[27] .is_wysiwyg = "true";
defparam \E_src2_imm[27] .power_up = "low";

cyclonev_lcell_comb \Add8~125 (
	.dataa(!\E_ctrl_alu_subtract~q ),
	.datab(!\E_ctrl_src2_choose_imm~q ),
	.datac(!\E_stw_data[27]~37_combout ),
	.datad(!\E_src2_imm[27]~q ),
	.datae(gnd),
	.dataf(!\E_src1[27]~55_combout ),
	.datag(gnd),
	.cin(\Add8~130 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add8~125_sumout ),
	.cout(\Add8~126 ),
	.shareout());
defparam \Add8~125 .extended_lut = "off";
defparam \Add8~125 .lut_mask = 64'h0000FF0000006996;
defparam \Add8~125 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_prelim[27]~28 (
	.dataa(!\M_wr_data_unfiltered[27]~25_combout ),
	.datab(!\D_src2_hazard_M~combout ),
	.datac(!\D_src2_hazard_W~combout ),
	.datad(!\W_wr_data[27]~q ),
	.datae(!\processor_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[27] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_prelim[27]~28_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_prelim[27]~28 .extended_lut = "off";
defparam \D_src2_prelim[27]~28 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \D_src2_prelim[27]~28 .shared_arith = "off";

dffeas \E_src2_prelim[27] (
	.clk(clk_clk),
	.d(\D_src2_prelim[27]~28_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_src2_prelim[27]~q ),
	.prn(vcc));
defparam \E_src2_prelim[27] .is_wysiwyg = "true";
defparam \E_src2_prelim[27] .power_up = "low";

cyclonev_lcell_comb \E_arith_src2[27]~18 (
	.dataa(!\E_src2_hazard_M~q ),
	.datab(!\E_ctrl_src2_choose_imm~q ),
	.datac(!\M_wr_data_unfiltered[27]~25_combout ),
	.datad(!\E_src2_imm[27]~q ),
	.datae(!\E_src2_prelim[27]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_arith_src2[27]~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_arith_src2[27]~18 .extended_lut = "off";
defparam \E_arith_src2[27]~18 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \E_arith_src2[27]~18 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[27]~50 (
	.dataa(!\E_compare_op[1]~q ),
	.datab(!\E_compare_op[0]~q ),
	.datac(!\E_arith_src2[27]~18_combout ),
	.datad(!\E_src1[27]~55_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[27]~50_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[27]~50 .extended_lut = "off";
defparam \E_alu_result[27]~50 .lut_mask = 64'h6996699669966996;
defparam \E_alu_result[27]~50 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[27]~51 (
	.dataa(!\E_ctrl_logic~q ),
	.datab(!\E_alu_result~0_combout ),
	.datac(!\Add8~125_sumout ),
	.datad(!\E_alu_result[27]~50_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[27]~51_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[27]~51 .extended_lut = "off";
defparam \E_alu_result[27]~51 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \E_alu_result[27]~51 .shared_arith = "off";

dffeas \M_alu_result[27] (
	.clk(clk_clk),
	.d(\E_alu_result[27]~51_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\M_alu_result[27]~q ),
	.prn(vcc));
defparam \M_alu_result[27] .is_wysiwyg = "true";
defparam \M_alu_result[27] .power_up = "low";

cyclonev_lcell_comb \M_wr_data_unfiltered[27]~25 (
	.dataa(!\M_ctrl_shift_rot~q ),
	.datab(!\av_ld_or_div_done~q ),
	.datac(!\M_shift_rot_result[27]~q ),
	.datad(!\av_ld_data_aligned_or_div[27]~q ),
	.datae(!\M_alu_result[27]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_wr_data_unfiltered[27]~25_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_wr_data_unfiltered[27]~25 .extended_lut = "off";
defparam \M_wr_data_unfiltered[27]~25 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \M_wr_data_unfiltered[27]~25 .shared_arith = "off";

cyclonev_lcell_comb \E_stw_data[27]~37 (
	.dataa(!\E_src2_hazard_M~q ),
	.datab(!\M_wr_data_unfiltered[27]~25_combout ),
	.datac(!\E_src2_prelim[27]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_stw_data[27]~37_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_stw_data[27]~37 .extended_lut = "off";
defparam \E_stw_data[27]~37 .lut_mask = 64'h2727272727272727;
defparam \E_stw_data[27]~37 .shared_arith = "off";

cyclonev_lcell_comb \Add8~101 (
	.dataa(!\E_ctrl_alu_subtract~q ),
	.datab(!\E_ctrl_src2_choose_imm~q ),
	.datac(!\E_stw_data[28]~28_combout ),
	.datad(!\E_src2_imm[28]~q ),
	.datae(gnd),
	.dataf(!\E_src1[28]~43_combout ),
	.datag(gnd),
	.cin(\Add8~126 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add8~101_sumout ),
	.cout(\Add8~102 ),
	.shareout());
defparam \Add8~101 .extended_lut = "off";
defparam \Add8~101 .lut_mask = 64'h0000FF0000006996;
defparam \Add8~101 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[28]~42 (
	.dataa(!\E_ctrl_src2_choose_imm~q ),
	.datab(!\E_compare_op[1]~q ),
	.datac(!\E_compare_op[0]~q ),
	.datad(!\E_src1[28]~43_combout ),
	.datae(!\E_src2_imm[28]~q ),
	.dataf(!\E_stw_data[28]~28_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[28]~42_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[28]~42 .extended_lut = "off";
defparam \E_alu_result[28]~42 .lut_mask = 64'h6996966996696996;
defparam \E_alu_result[28]~42 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[28]~43 (
	.dataa(!\E_ctrl_logic~q ),
	.datab(!\E_alu_result~0_combout ),
	.datac(!\Add8~101_sumout ),
	.datad(!\E_alu_result[28]~42_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[28]~43_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[28]~43 .extended_lut = "off";
defparam \E_alu_result[28]~43 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \E_alu_result[28]~43 .shared_arith = "off";

dffeas \M_alu_result[28] (
	.clk(clk_clk),
	.d(\E_alu_result[28]~43_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\M_alu_result[28]~q ),
	.prn(vcc));
defparam \M_alu_result[28] .is_wysiwyg = "true";
defparam \M_alu_result[28] .power_up = "low";

cyclonev_lcell_comb \E_src1[28]~41 (
	.dataa(!\M_ctrl_shift_rot~q ),
	.datab(!\av_ld_or_div_done~q ),
	.datac(!\E_src1_hazard_M~q ),
	.datad(!\M_shift_rot_result[28]~q ),
	.datae(!\av_ld_data_aligned_or_div[28]~q ),
	.dataf(!\M_alu_result[28]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_src1[28]~41_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_src1[28]~41 .extended_lut = "off";
defparam \E_src1[28]~41 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \E_src1[28]~41 .shared_arith = "off";

cyclonev_lcell_comb \D_src1_prelim[28]~23 (
	.dataa(!\M_wr_data_unfiltered[28]~29_combout ),
	.datab(!\D_src1_hazard_M~combout ),
	.datac(!\D_src1_hazard_W~combout ),
	.datad(!\W_wr_data[28]~q ),
	.datae(!\processor_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[28] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_prelim[28]~23_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src1_prelim[28]~23 .extended_lut = "off";
defparam \D_src1_prelim[28]~23 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \D_src1_prelim[28]~23 .shared_arith = "off";

dffeas \E_src1_prelim[28] (
	.clk(clk_clk),
	.d(\D_src1_prelim[28]~23_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_src1_prelim[28]~q ),
	.prn(vcc));
defparam \E_src1_prelim[28] .is_wysiwyg = "true";
defparam \E_src1_prelim[28] .power_up = "low";

cyclonev_lcell_comb \E_src1[28]~42 (
	.dataa(!\E_src1_hazard_M~q ),
	.datab(!\E_src1_prelim[28]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_src1[28]~42_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_src1[28]~42 .extended_lut = "off";
defparam \E_src1[28]~42 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \E_src1[28]~42 .shared_arith = "off";

cyclonev_lcell_comb \E_src1[28]~43 (
	.dataa(!\E_src1[28]~41_combout ),
	.datab(!\E_src1[28]~42_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_src1[28]~43_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_src1[28]~43 .extended_lut = "off";
defparam \E_src1[28]~43 .lut_mask = 64'h7777777777777777;
defparam \E_src1[28]~43 .shared_arith = "off";

cyclonev_lcell_comb \M_shift_rot_result_nxt[28]~23 (
	.dataa(!\M_shift_rot_stall~q ),
	.datab(!\M_ctrl_shift_rot_right~q ),
	.datac(!\M_shift_rot_result[29]~q ),
	.datad(!\E_src1[28]~43_combout ),
	.datae(!\M_shift_rot_result[27]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_shift_rot_result_nxt[28]~23_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_shift_rot_result_nxt[28]~23 .extended_lut = "off";
defparam \M_shift_rot_result_nxt[28]~23 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \M_shift_rot_result_nxt[28]~23 .shared_arith = "off";

dffeas \M_shift_rot_result[28] (
	.clk(clk_clk),
	.d(\M_shift_rot_result_nxt[28]~23_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\M_shift_rot_result[28]~q ),
	.prn(vcc));
defparam \M_shift_rot_result[28] .is_wysiwyg = "true";
defparam \M_shift_rot_result[28] .power_up = "low";

dffeas \W_wr_data[29] (
	.clk(clk_clk),
	.d(\M_wr_data_unfiltered[29]~20_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\W_wr_data[29]~q ),
	.prn(vcc));
defparam \W_wr_data[29] .is_wysiwyg = "true";
defparam \W_wr_data[29] .power_up = "low";

cyclonev_lcell_comb \D_src1_prelim[29]~21 (
	.dataa(!\M_wr_data_unfiltered[29]~20_combout ),
	.datab(!\D_src1_hazard_M~combout ),
	.datac(!\D_src1_hazard_W~combout ),
	.datad(!\W_wr_data[29]~q ),
	.datae(!\processor_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[29] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_prelim[29]~21_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src1_prelim[29]~21 .extended_lut = "off";
defparam \D_src1_prelim[29]~21 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \D_src1_prelim[29]~21 .shared_arith = "off";

dffeas \E_src1_prelim[29] (
	.clk(clk_clk),
	.d(\D_src1_prelim[29]~21_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_src1_prelim[29]~q ),
	.prn(vcc));
defparam \E_src1_prelim[29] .is_wysiwyg = "true";
defparam \E_src1_prelim[29] .power_up = "low";

cyclonev_lcell_comb \E_src1[29]~39 (
	.dataa(!\E_src1_hazard_M~q ),
	.datab(!\M_wr_data_unfiltered[29]~20_combout ),
	.datac(!\E_src1_prelim[29]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_src1[29]~39_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_src1[29]~39 .extended_lut = "off";
defparam \E_src1[29]~39 .lut_mask = 64'h2727272727272727;
defparam \E_src1[29]~39 .shared_arith = "off";

cyclonev_lcell_comb \M_shift_rot_result_nxt[29]~21 (
	.dataa(!\M_shift_rot_stall~q ),
	.datab(!\M_ctrl_shift_rot_right~q ),
	.datac(!\M_shift_rot_result[30]~q ),
	.datad(!\M_shift_rot_result[28]~q ),
	.datae(!\E_src1[29]~39_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_shift_rot_result_nxt[29]~21_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_shift_rot_result_nxt[29]~21 .extended_lut = "off";
defparam \M_shift_rot_result_nxt[29]~21 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \M_shift_rot_result_nxt[29]~21 .shared_arith = "off";

dffeas \M_shift_rot_result[29] (
	.clk(clk_clk),
	.d(\M_shift_rot_result_nxt[29]~21_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\M_shift_rot_result[29]~q ),
	.prn(vcc));
defparam \M_shift_rot_result[29] .is_wysiwyg = "true";
defparam \M_shift_rot_result[29] .power_up = "low";

dffeas \av_ld_data_aligned_or_div[29] (
	.clk(clk_clk),
	.d(\av_fill_bit~0_combout ),
	.asdata(\d_readdata_d1[29]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\M_iw[4]~q ),
	.ena(vcc),
	.q(\av_ld_data_aligned_or_div[29]~q ),
	.prn(vcc));
defparam \av_ld_data_aligned_or_div[29] .is_wysiwyg = "true";
defparam \av_ld_data_aligned_or_div[29] .power_up = "low";

dffeas \E_src2_imm[29] (
	.clk(clk_clk),
	.d(\D_iw[21]~q ),
	.asdata(\D_iw[19]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\D_ctrl_unsigned_lo_imm16~combout ),
	.sload(\Equal171~0_combout ),
	.ena(\W_stall~combout ),
	.q(\E_src2_imm[29]~q ),
	.prn(vcc));
defparam \E_src2_imm[29] .is_wysiwyg = "true";
defparam \E_src2_imm[29] .power_up = "low";

cyclonev_lcell_comb \Add8~89 (
	.dataa(!\E_ctrl_alu_subtract~q ),
	.datab(!\E_ctrl_src2_choose_imm~q ),
	.datac(!\E_stw_data[29]~22_combout ),
	.datad(!\E_src2_imm[29]~q ),
	.datae(gnd),
	.dataf(!\E_src1[29]~39_combout ),
	.datag(gnd),
	.cin(\Add8~102 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add8~89_sumout ),
	.cout(\Add8~90 ),
	.shareout());
defparam \Add8~89 .extended_lut = "off";
defparam \Add8~89 .lut_mask = 64'h0000FF0000006996;
defparam \Add8~89 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_prelim[29]~22 (
	.dataa(!\M_wr_data_unfiltered[29]~20_combout ),
	.datab(!\D_src2_hazard_M~combout ),
	.datac(!\D_src2_hazard_W~combout ),
	.datad(!\W_wr_data[29]~q ),
	.datae(!\processor_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[29] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_prelim[29]~22_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_prelim[29]~22 .extended_lut = "off";
defparam \D_src2_prelim[29]~22 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \D_src2_prelim[29]~22 .shared_arith = "off";

dffeas \E_src2_prelim[29] (
	.clk(clk_clk),
	.d(\D_src2_prelim[29]~22_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_src2_prelim[29]~q ),
	.prn(vcc));
defparam \E_src2_prelim[29] .is_wysiwyg = "true";
defparam \E_src2_prelim[29] .power_up = "low";

cyclonev_lcell_comb \E_arith_src2[29]~14 (
	.dataa(!\E_src2_hazard_M~q ),
	.datab(!\E_ctrl_src2_choose_imm~q ),
	.datac(!\M_wr_data_unfiltered[29]~20_combout ),
	.datad(!\E_src2_imm[29]~q ),
	.datae(!\E_src2_prelim[29]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_arith_src2[29]~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_arith_src2[29]~14 .extended_lut = "off";
defparam \E_arith_src2[29]~14 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \E_arith_src2[29]~14 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[29]~34 (
	.dataa(!\E_compare_op[1]~q ),
	.datab(!\E_compare_op[0]~q ),
	.datac(!\E_arith_src2[29]~14_combout ),
	.datad(!\E_src1[29]~39_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[29]~34_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[29]~34 .extended_lut = "off";
defparam \E_alu_result[29]~34 .lut_mask = 64'h6996699669966996;
defparam \E_alu_result[29]~34 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[29]~35 (
	.dataa(!\E_ctrl_logic~q ),
	.datab(!\E_alu_result~0_combout ),
	.datac(!\Add8~89_sumout ),
	.datad(!\E_alu_result[29]~34_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[29]~35_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[29]~35 .extended_lut = "off";
defparam \E_alu_result[29]~35 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \E_alu_result[29]~35 .shared_arith = "off";

dffeas \M_alu_result[29] (
	.clk(clk_clk),
	.d(\E_alu_result[29]~35_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\M_alu_result[29]~q ),
	.prn(vcc));
defparam \M_alu_result[29] .is_wysiwyg = "true";
defparam \M_alu_result[29] .power_up = "low";

cyclonev_lcell_comb \M_wr_data_unfiltered[29]~20 (
	.dataa(!\M_ctrl_shift_rot~q ),
	.datab(!\av_ld_or_div_done~q ),
	.datac(!\M_shift_rot_result[29]~q ),
	.datad(!\av_ld_data_aligned_or_div[29]~q ),
	.datae(!\M_alu_result[29]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_wr_data_unfiltered[29]~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_wr_data_unfiltered[29]~20 .extended_lut = "off";
defparam \M_wr_data_unfiltered[29]~20 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \M_wr_data_unfiltered[29]~20 .shared_arith = "off";

cyclonev_lcell_comb \E_stw_data[29]~22 (
	.dataa(!\E_src2_hazard_M~q ),
	.datab(!\M_wr_data_unfiltered[29]~20_combout ),
	.datac(!\E_src2_prelim[29]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_stw_data[29]~22_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_stw_data[29]~22 .extended_lut = "off";
defparam \E_stw_data[29]~22 .lut_mask = 64'h2727272727272727;
defparam \E_stw_data[29]~22 .shared_arith = "off";

cyclonev_lcell_comb \Add8~81 (
	.dataa(!\E_ctrl_alu_subtract~q ),
	.datab(!\E_ctrl_src2_choose_imm~q ),
	.datac(!\E_stw_data[30]~17_combout ),
	.datad(!\E_src2_imm[30]~q ),
	.datae(gnd),
	.dataf(!\E_src1[30]~35_combout ),
	.datag(gnd),
	.cin(\Add8~90 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add8~81_sumout ),
	.cout(\Add8~82 ),
	.shareout());
defparam \Add8~81 .extended_lut = "off";
defparam \Add8~81 .lut_mask = 64'h0000FF0000006996;
defparam \Add8~81 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[30]~30 (
	.dataa(!\E_ctrl_src2_choose_imm~q ),
	.datab(!\E_compare_op[1]~q ),
	.datac(!\E_compare_op[0]~q ),
	.datad(!\E_src1[30]~35_combout ),
	.datae(!\E_src2_imm[30]~q ),
	.dataf(!\E_stw_data[30]~17_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[30]~30_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[30]~30 .extended_lut = "off";
defparam \E_alu_result[30]~30 .lut_mask = 64'h6996966996696996;
defparam \E_alu_result[30]~30 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[30]~31 (
	.dataa(!\E_ctrl_logic~q ),
	.datab(!\E_alu_result~0_combout ),
	.datac(!\Add8~81_sumout ),
	.datad(!\E_alu_result[30]~30_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[30]~31_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[30]~31 .extended_lut = "off";
defparam \E_alu_result[30]~31 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \E_alu_result[30]~31 .shared_arith = "off";

dffeas \M_alu_result[30] (
	.clk(clk_clk),
	.d(\E_alu_result[30]~31_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\M_alu_result[30]~q ),
	.prn(vcc));
defparam \M_alu_result[30] .is_wysiwyg = "true";
defparam \M_alu_result[30] .power_up = "low";

cyclonev_lcell_comb \E_src1[30]~33 (
	.dataa(!\M_ctrl_shift_rot~q ),
	.datab(!\av_ld_or_div_done~q ),
	.datac(!\E_src1_hazard_M~q ),
	.datad(!\M_shift_rot_result[30]~q ),
	.datae(!\av_ld_data_aligned_or_div[30]~q ),
	.dataf(!\M_alu_result[30]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_src1[30]~33_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_src1[30]~33 .extended_lut = "off";
defparam \E_src1[30]~33 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \E_src1[30]~33 .shared_arith = "off";

cyclonev_lcell_comb \D_src1_prelim[30]~19 (
	.dataa(!\M_wr_data_unfiltered[30]~19_combout ),
	.datab(!\D_src1_hazard_M~combout ),
	.datac(!\D_src1_hazard_W~combout ),
	.datad(!\W_wr_data[30]~q ),
	.datae(!\processor_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[30] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_prelim[30]~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src1_prelim[30]~19 .extended_lut = "off";
defparam \D_src1_prelim[30]~19 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \D_src1_prelim[30]~19 .shared_arith = "off";

dffeas \E_src1_prelim[30] (
	.clk(clk_clk),
	.d(\D_src1_prelim[30]~19_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_src1_prelim[30]~q ),
	.prn(vcc));
defparam \E_src1_prelim[30] .is_wysiwyg = "true";
defparam \E_src1_prelim[30] .power_up = "low";

cyclonev_lcell_comb \E_src1[30]~34 (
	.dataa(!\E_src1_hazard_M~q ),
	.datab(!\E_src1_prelim[30]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_src1[30]~34_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_src1[30]~34 .extended_lut = "off";
defparam \E_src1[30]~34 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \E_src1[30]~34 .shared_arith = "off";

cyclonev_lcell_comb \E_src1[30]~35 (
	.dataa(!\E_src1[30]~33_combout ),
	.datab(!\E_src1[30]~34_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_src1[30]~35_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_src1[30]~35 .extended_lut = "off";
defparam \E_src1[30]~35 .lut_mask = 64'h7777777777777777;
defparam \E_src1[30]~35 .shared_arith = "off";

cyclonev_lcell_comb \M_shift_rot_result_nxt[30]~19 (
	.dataa(!\M_shift_rot_stall~q ),
	.datab(!\M_ctrl_shift_rot_right~q ),
	.datac(!\M_shift_rot_result[31]~q ),
	.datad(!\E_src1[30]~35_combout ),
	.datae(!\M_shift_rot_result[29]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_shift_rot_result_nxt[30]~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_shift_rot_result_nxt[30]~19 .extended_lut = "off";
defparam \M_shift_rot_result_nxt[30]~19 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \M_shift_rot_result_nxt[30]~19 .shared_arith = "off";

dffeas \M_shift_rot_result[30] (
	.clk(clk_clk),
	.d(\M_shift_rot_result_nxt[30]~19_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\M_shift_rot_result[30]~q ),
	.prn(vcc));
defparam \M_shift_rot_result[30] .is_wysiwyg = "true";
defparam \M_shift_rot_result[30] .power_up = "low";

dffeas \W_wr_data[31] (
	.clk(clk_clk),
	.d(\M_wr_data_unfiltered[31]~17_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\W_wr_data[31]~q ),
	.prn(vcc));
defparam \W_wr_data[31] .is_wysiwyg = "true";
defparam \W_wr_data[31] .power_up = "low";

cyclonev_lcell_comb \D_src1_prelim[31]~17 (
	.dataa(!\M_wr_data_unfiltered[31]~17_combout ),
	.datab(!\D_src1_hazard_M~combout ),
	.datac(!\D_src1_hazard_W~combout ),
	.datad(!\W_wr_data[31]~q ),
	.datae(!\processor_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[31] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_prelim[31]~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src1_prelim[31]~17 .extended_lut = "off";
defparam \D_src1_prelim[31]~17 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \D_src1_prelim[31]~17 .shared_arith = "off";

dffeas \E_src1_prelim[31] (
	.clk(clk_clk),
	.d(\D_src1_prelim[31]~17_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_src1_prelim[31]~q ),
	.prn(vcc));
defparam \E_src1_prelim[31] .is_wysiwyg = "true";
defparam \E_src1_prelim[31] .power_up = "low";

cyclonev_lcell_comb \E_src1[31]~31 (
	.dataa(!\E_src1_hazard_M~q ),
	.datab(!\M_wr_data_unfiltered[31]~17_combout ),
	.datac(!\E_src1_prelim[31]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_src1[31]~31_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_src1[31]~31 .extended_lut = "off";
defparam \E_src1[31]~31 .lut_mask = 64'h2727272727272727;
defparam \E_src1[31]~31 .shared_arith = "off";

cyclonev_lcell_comb \M_shift_rot_result_nxt[31]~17 (
	.dataa(!\M_shift_rot_stall~q ),
	.datab(!\M_ctrl_shift_rot_right~q ),
	.datac(!\M_shift_rot_fill_bit~0_combout ),
	.datad(!\M_shift_rot_result[30]~q ),
	.datae(!\E_src1[31]~31_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_shift_rot_result_nxt[31]~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_shift_rot_result_nxt[31]~17 .extended_lut = "off";
defparam \M_shift_rot_result_nxt[31]~17 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \M_shift_rot_result_nxt[31]~17 .shared_arith = "off";

dffeas \M_shift_rot_result[31] (
	.clk(clk_clk),
	.d(\M_shift_rot_result_nxt[31]~17_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\M_shift_rot_result[31]~q ),
	.prn(vcc));
defparam \M_shift_rot_result[31] .is_wysiwyg = "true";
defparam \M_shift_rot_result[31] .power_up = "low";

dffeas \av_ld_data_aligned_or_div[31] (
	.clk(clk_clk),
	.d(\av_fill_bit~0_combout ),
	.asdata(\d_readdata_d1[31]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\M_iw[4]~q ),
	.ena(vcc),
	.q(\av_ld_data_aligned_or_div[31]~q ),
	.prn(vcc));
defparam \av_ld_data_aligned_or_div[31] .is_wysiwyg = "true";
defparam \av_ld_data_aligned_or_div[31] .power_up = "low";

cyclonev_lcell_comb \Equal4~14 (
	.dataa(!\D_iw[0]~q ),
	.datab(!\D_iw[1]~q ),
	.datac(!\D_iw[2]~q ),
	.datad(!\D_iw[3]~q ),
	.datae(!\D_iw[4]~q ),
	.dataf(!\D_iw[5]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal4~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal4~14 .extended_lut = "off";
defparam \Equal4~14 .lut_mask = 64'hFFFFFFFFFFFFBFFF;
defparam \Equal4~14 .shared_arith = "off";

cyclonev_lcell_comb \Equal4~15 (
	.dataa(!\D_iw[0]~q ),
	.datab(!\D_iw[1]~q ),
	.datac(!\D_iw[2]~q ),
	.datad(!\D_iw[3]~q ),
	.datae(!\D_iw[4]~q ),
	.dataf(!\D_iw[5]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal4~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal4~15 .extended_lut = "off";
defparam \Equal4~15 .lut_mask = 64'hFFFFFFFFFFBFFFFF;
defparam \Equal4~15 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_alu_signed_comparison~0 (
	.dataa(!\D_iw[16]~q ),
	.datab(!\D_iw[15]~q ),
	.datac(!\D_iw[14]~q ),
	.datad(!\D_iw[11]~q ),
	.datae(!\D_ctrl_cmp~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_alu_signed_comparison~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_alu_signed_comparison~0 .extended_lut = "off";
defparam \D_ctrl_alu_signed_comparison~0 .lut_mask = 64'hFFBEFFFFFFBEFFFF;
defparam \D_ctrl_alu_signed_comparison~0 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_alu_signed_comparison~1 (
	.dataa(!\Equal4~9_combout ),
	.datab(!\Equal4~10_combout ),
	.datac(!\Equal4~14_combout ),
	.datad(!\Equal4~15_combout ),
	.datae(!\D_ctrl_alu_signed_comparison~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_alu_signed_comparison~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_alu_signed_comparison~1 .extended_lut = "off";
defparam \D_ctrl_alu_signed_comparison~1 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \D_ctrl_alu_signed_comparison~1 .shared_arith = "off";

dffeas E_ctrl_alu_signed_comparison(
	.clk(clk_clk),
	.d(\D_ctrl_alu_signed_comparison~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_ctrl_alu_signed_comparison~q ),
	.prn(vcc));
defparam E_ctrl_alu_signed_comparison.is_wysiwyg = "true";
defparam E_ctrl_alu_signed_comparison.power_up = "low";

cyclonev_lcell_comb \D_src2_imm[31]~0 (
	.dataa(!\D_iw[21]~q ),
	.datab(!\D_ctrl_unsigned_lo_imm16~combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_imm[31]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_imm[31]~0 .extended_lut = "off";
defparam \D_src2_imm[31]~0 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \D_src2_imm[31]~0 .shared_arith = "off";

dffeas \E_src2_imm[31] (
	.clk(clk_clk),
	.d(\D_src2_imm[31]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_src2_imm[31]~q ),
	.prn(vcc));
defparam \E_src2_imm[31] .is_wysiwyg = "true";
defparam \E_src2_imm[31] .power_up = "low";

cyclonev_lcell_comb \D_src2_prelim[31]~17 (
	.dataa(!\M_wr_data_unfiltered[31]~17_combout ),
	.datab(!\D_src2_hazard_M~combout ),
	.datac(!\D_src2_hazard_W~combout ),
	.datad(!\W_wr_data[31]~q ),
	.datae(!\processor_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[31] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_prelim[31]~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_prelim[31]~17 .extended_lut = "off";
defparam \D_src2_prelim[31]~17 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \D_src2_prelim[31]~17 .shared_arith = "off";

dffeas \E_src2_prelim[31] (
	.clk(clk_clk),
	.d(\D_src2_prelim[31]~17_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_src2_prelim[31]~q ),
	.prn(vcc));
defparam \E_src2_prelim[31] .is_wysiwyg = "true";
defparam \E_src2_prelim[31] .power_up = "low";

cyclonev_lcell_comb \E_src2[31]~0 (
	.dataa(!\E_src2_hazard_M~q ),
	.datab(!\E_ctrl_src2_choose_imm~q ),
	.datac(!\M_wr_data_unfiltered[31]~17_combout ),
	.datad(!\E_src2_imm[31]~q ),
	.datae(!\E_src2_prelim[31]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_src2[31]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_src2[31]~0 .extended_lut = "off";
defparam \E_src2[31]~0 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \E_src2[31]~0 .shared_arith = "off";

cyclonev_lcell_comb \Add8~73 (
	.dataa(!\E_ctrl_alu_signed_comparison~q ),
	.datab(!\E_ctrl_alu_subtract~q ),
	.datac(gnd),
	.datad(!\E_src2[31]~0_combout ),
	.datae(gnd),
	.dataf(!\E_src1[31]~31_combout ),
	.datag(gnd),
	.cin(\Add8~82 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add8~73_sumout ),
	.cout(\Add8~74 ),
	.shareout());
defparam \Add8~73 .extended_lut = "off";
defparam \Add8~73 .lut_mask = 64'h000055AA00009966;
defparam \Add8~73 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[31]~26 (
	.dataa(!\E_compare_op[1]~q ),
	.datab(!\E_compare_op[0]~q ),
	.datac(!\E_src2[31]~0_combout ),
	.datad(!\E_src1[31]~31_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[31]~26_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[31]~26 .extended_lut = "off";
defparam \E_alu_result[31]~26 .lut_mask = 64'h6996699669966996;
defparam \E_alu_result[31]~26 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[31]~27 (
	.dataa(!\E_ctrl_logic~q ),
	.datab(!\E_alu_result~0_combout ),
	.datac(!\Add8~73_sumout ),
	.datad(!\E_alu_result[31]~26_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[31]~27_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[31]~27 .extended_lut = "off";
defparam \E_alu_result[31]~27 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \E_alu_result[31]~27 .shared_arith = "off";

dffeas \M_alu_result[31] (
	.clk(clk_clk),
	.d(\E_alu_result[31]~27_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\M_alu_result[31]~q ),
	.prn(vcc));
defparam \M_alu_result[31] .is_wysiwyg = "true";
defparam \M_alu_result[31] .power_up = "low";

cyclonev_lcell_comb \M_wr_data_unfiltered[31]~17 (
	.dataa(!\M_ctrl_shift_rot~q ),
	.datab(!\av_ld_or_div_done~q ),
	.datac(!\M_shift_rot_result[31]~q ),
	.datad(!\av_ld_data_aligned_or_div[31]~q ),
	.datae(!\M_alu_result[31]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_wr_data_unfiltered[31]~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_wr_data_unfiltered[31]~17 .extended_lut = "off";
defparam \M_wr_data_unfiltered[31]~17 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \M_wr_data_unfiltered[31]~17 .shared_arith = "off";

cyclonev_lcell_comb \E_logic_result~0 (
	.dataa(!\E_ctrl_src2_choose_imm~q ),
	.datab(!\E_src1[30]~33_combout ),
	.datac(!\E_src1[30]~34_combout ),
	.datad(!\E_src2_imm[30]~q ),
	.datae(!\E_stw_data[30]~15_combout ),
	.dataf(!\E_stw_data[30]~16_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_logic_result~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_logic_result~0 .extended_lut = "off";
defparam \E_logic_result~0 .lut_mask = 64'h6996966996696996;
defparam \E_logic_result~0 .shared_arith = "off";

cyclonev_lcell_comb \E_logic_result~1 (
	.dataa(!\E_ctrl_src2_choose_imm~q ),
	.datab(!\E_src1[28]~41_combout ),
	.datac(!\E_src1[28]~42_combout ),
	.datad(!\E_src2_imm[28]~q ),
	.datae(!\E_stw_data[28]~26_combout ),
	.dataf(!\E_stw_data[28]~27_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_logic_result~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_logic_result~1 .extended_lut = "off";
defparam \E_logic_result~1 .lut_mask = 64'h6996966996696996;
defparam \E_logic_result~1 .shared_arith = "off";

cyclonev_lcell_comb \E_logic_result~2 (
	.dataa(!\E_ctrl_src2_choose_imm~q ),
	.datab(!\E_src1[26]~56_combout ),
	.datac(!\E_src1[26]~57_combout ),
	.datad(!\E_src2_imm[26]~q ),
	.datae(!\E_stw_data[26]~38_combout ),
	.dataf(!\E_stw_data[26]~39_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_logic_result~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_logic_result~2 .extended_lut = "off";
defparam \E_logic_result~2 .lut_mask = 64'h6996966996696996;
defparam \E_logic_result~2 .shared_arith = "off";

cyclonev_lcell_comb \E_logic_result~3 (
	.dataa(!\E_ctrl_src2_choose_imm~q ),
	.datab(!\E_src1[24]~44_combout ),
	.datac(!\E_src1[24]~45_combout ),
	.datad(!\E_src2_imm[24]~q ),
	.datae(!\E_stw_data[24]~18_combout ),
	.dataf(!\E_stw_data[24]~19_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_logic_result~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_logic_result~3 .extended_lut = "off";
defparam \E_logic_result~3 .lut_mask = 64'h6996966996696996;
defparam \E_logic_result~3 .shared_arith = "off";

cyclonev_lcell_comb \E_logic_result~4 (
	.dataa(!\E_ctrl_src2_choose_imm~q ),
	.datab(!\E_src1[22]~51_combout ),
	.datac(!\E_src1[22]~52_combout ),
	.datad(!\E_src2_imm[22]~q ),
	.datae(!\E_stw_data[22]~29_combout ),
	.dataf(!\E_stw_data[22]~30_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_logic_result~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_logic_result~4 .extended_lut = "off";
defparam \E_logic_result~4 .lut_mask = 64'h6996966996696996;
defparam \E_logic_result~4 .shared_arith = "off";

cyclonev_lcell_comb \E_logic_result~5 (
	.dataa(!\E_ctrl_src2_choose_imm~q ),
	.datab(!\E_src1[20]~48_combout ),
	.datac(!\E_src1[20]~49_combout ),
	.datad(!\E_src2_imm[20]~q ),
	.datae(!\E_stw_data[20]~23_combout ),
	.dataf(!\E_stw_data[20]~24_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_logic_result~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_logic_result~5 .extended_lut = "off";
defparam \E_logic_result~5 .lut_mask = 64'h6996966996696996;
defparam \E_logic_result~5 .shared_arith = "off";

cyclonev_lcell_comb \E_logic_result~6 (
	.dataa(!\E_ctrl_src2_choose_imm~q ),
	.datab(!\E_src1[18]~36_combout ),
	.datac(!\E_src1[18]~37_combout ),
	.datad(!\E_src2_imm[18]~q ),
	.datae(!\E_stw_data[18]~32_combout ),
	.dataf(!\E_stw_data[18]~33_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_logic_result~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_logic_result~6 .extended_lut = "off";
defparam \E_logic_result~6 .lut_mask = 64'h6996966996696996;
defparam \E_logic_result~6 .shared_arith = "off";

cyclonev_lcell_comb \E_logic_result~7 (
	.dataa(!\E_ctrl_src2_choose_imm~q ),
	.datab(!\E_stw_data[16]~0_combout ),
	.datac(!\E_stw_data[16]~1_combout ),
	.datad(!\E_src2_imm[16]~q ),
	.datae(!\E_src1[16]~7_combout ),
	.dataf(!\E_src1[16]~8_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_logic_result~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_logic_result~7 .extended_lut = "off";
defparam \E_logic_result~7 .lut_mask = 64'h6996966996696996;
defparam \E_logic_result~7 .shared_arith = "off";

cyclonev_lcell_comb \E_arith_src2[15]~2 (
	.dataa(!\E_ctrl_src2_choose_imm~q ),
	.datab(!\E_src2_imm[15]~q ),
	.datac(!\E_src2_hazard_M~q ),
	.datad(!\M_wr_data_unfiltered[15]~1_combout ),
	.datae(!\E_src2_prelim[15]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_arith_src2[15]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_arith_src2[15]~2 .extended_lut = "off";
defparam \E_arith_src2[15]~2 .lut_mask = 64'h7BFFFFFF7BFFFFFF;
defparam \E_arith_src2[15]~2 .shared_arith = "off";

cyclonev_lcell_comb \E_logic_result~18 (
	.dataa(!\E_src1_prelim[14]~q ),
	.datab(!\E_src2_prelim[14]~q ),
	.datac(!\E_src2_imm[14]~q ),
	.datad(!\E_src1_hazard_M~q ),
	.datae(!\E_ctrl_src2_choose_imm~q ),
	.dataf(!\M_wr_data_unfiltered[14]~2_combout ),
	.datag(!\E_src2_hazard_M~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_logic_result~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_logic_result~18 .extended_lut = "on";
defparam \E_logic_result~18 .lut_mask = 64'h6996699669966996;
defparam \E_logic_result~18 .shared_arith = "off";

cyclonev_lcell_comb \E_arith_src2[13]~4 (
	.dataa(!\E_src2_hazard_M~q ),
	.datab(!\E_ctrl_src2_choose_imm~q ),
	.datac(!\M_wr_data_unfiltered[13]~3_combout ),
	.datad(!\E_src2_prelim[13]~q ),
	.datae(!\E_src2_imm[13]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_arith_src2[13]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_arith_src2[13]~4 .extended_lut = "off";
defparam \E_arith_src2[13]~4 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \E_arith_src2[13]~4 .shared_arith = "off";

cyclonev_lcell_comb \E_logic_result~14 (
	.dataa(!\E_src1_prelim[12]~q ),
	.datab(!\E_src2_prelim[12]~q ),
	.datac(!\E_src2_imm[12]~q ),
	.datad(!\E_src1_hazard_M~q ),
	.datae(!\E_ctrl_src2_choose_imm~q ),
	.dataf(!\M_wr_data_unfiltered[12]~4_combout ),
	.datag(!\E_src2_hazard_M~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_logic_result~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_logic_result~14 .extended_lut = "on";
defparam \E_logic_result~14 .lut_mask = 64'h6996699669966996;
defparam \E_logic_result~14 .shared_arith = "off";

cyclonev_lcell_comb \E_arith_src2[11]~6 (
	.dataa(!\E_src2_hazard_M~q ),
	.datab(!\E_ctrl_src2_choose_imm~q ),
	.datac(!\M_wr_data_unfiltered[11]~5_combout ),
	.datad(!\E_src2_prelim[11]~q ),
	.datae(!\E_src2_imm[11]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_arith_src2[11]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_arith_src2[11]~6 .extended_lut = "off";
defparam \E_arith_src2[11]~6 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \E_arith_src2[11]~6 .shared_arith = "off";

cyclonev_lcell_comb \E_logic_result~8 (
	.dataa(!\E_ctrl_src2_choose_imm~q ),
	.datab(!\E_stw_data[10]~6_combout ),
	.datac(!\E_stw_data[10]~7_combout ),
	.datad(!\E_src2_imm[10]~q ),
	.datae(!\E_src1[10]~15_combout ),
	.dataf(!\E_src1[10]~16_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_logic_result~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_logic_result~8 .extended_lut = "off";
defparam \E_logic_result~8 .lut_mask = 64'h6996966996696996;
defparam \E_logic_result~8 .shared_arith = "off";

cyclonev_lcell_comb \E_arith_src2[9]~7 (
	.dataa(!\E_src2_hazard_M~q ),
	.datab(!\E_ctrl_src2_choose_imm~q ),
	.datac(!\M_wr_data_unfiltered[9]~6_combout ),
	.datad(!\E_src2_prelim[9]~q ),
	.datae(!\E_src2_imm[9]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_arith_src2[9]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_arith_src2[9]~7 .extended_lut = "off";
defparam \E_arith_src2[9]~7 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \E_arith_src2[9]~7 .shared_arith = "off";

cyclonev_lcell_comb \E_logic_result~9 (
	.dataa(!\E_ctrl_src2_choose_imm~q ),
	.datab(!\E_stw_data[8]~9_combout ),
	.datac(!\E_stw_data[8]~10_combout ),
	.datad(!\E_src2_imm[8]~q ),
	.datae(!\E_src1[8]~19_combout ),
	.dataf(!\E_src1[8]~20_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_logic_result~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_logic_result~9 .extended_lut = "off";
defparam \E_logic_result~9 .lut_mask = 64'h6996966996696996;
defparam \E_logic_result~9 .shared_arith = "off";

cyclonev_lcell_comb \E_arith_src2[7]~8 (
	.dataa(!\E_src2_hazard_M~q ),
	.datab(!\E_ctrl_src2_choose_imm~q ),
	.datac(!\M_wr_data_unfiltered[7]~7_combout ),
	.datad(!\E_src2_prelim[7]~q ),
	.datae(!\E_src2_imm[7]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_arith_src2[7]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_arith_src2[7]~8 .extended_lut = "off";
defparam \E_arith_src2[7]~8 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \E_arith_src2[7]~8 .shared_arith = "off";

cyclonev_lcell_comb \E_logic_result~10 (
	.dataa(!\E_ctrl_src2_choose_imm~q ),
	.datab(!\E_stb_data[6]~6_combout ),
	.datac(!\E_stb_data[6]~7_combout ),
	.datad(!\E_src2_imm[6]~q ),
	.datae(!\E_src1[6]~4_combout ),
	.dataf(!\E_src1[6]~5_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_logic_result~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_logic_result~10 .extended_lut = "off";
defparam \E_logic_result~10 .lut_mask = 64'h6996966996696996;
defparam \E_logic_result~10 .shared_arith = "off";

cyclonev_lcell_comb \E_arith_src2[5]~0 (
	.dataa(!\E_src2_hazard_M~q ),
	.datab(!\E_ctrl_src2_choose_imm~q ),
	.datac(!\M_wr_data_unfiltered[5]~0_combout ),
	.datad(!\E_src2_prelim[5]~q ),
	.datae(!\E_src2_imm[5]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_arith_src2[5]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_arith_src2[5]~0 .extended_lut = "off";
defparam \E_arith_src2[5]~0 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \E_arith_src2[5]~0 .shared_arith = "off";

cyclonev_lcell_comb \E_logic_result~11 (
	.dataa(!\E_ctrl_src2_choose_imm~q ),
	.datab(!\E_stb_data[4]~3_combout ),
	.datac(!\E_stb_data[4]~4_combout ),
	.datad(!\E_src2_imm[4]~q ),
	.datae(!\E_src1[4]~1_combout ),
	.dataf(!\E_src1[4]~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_logic_result~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_logic_result~11 .extended_lut = "off";
defparam \E_logic_result~11 .lut_mask = 64'h6996966996696996;
defparam \E_logic_result~11 .shared_arith = "off";

cyclonev_lcell_comb \E_arith_src2[3]~9 (
	.dataa(!\E_src2_hazard_M~q ),
	.datab(!\E_ctrl_src2_choose_imm~q ),
	.datac(!\M_wr_data_unfiltered[3]~8_combout ),
	.datad(!\E_src2_prelim[3]~q ),
	.datae(!\E_src2_imm[3]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_arith_src2[3]~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_arith_src2[3]~9 .extended_lut = "off";
defparam \E_arith_src2[3]~9 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \E_arith_src2[3]~9 .shared_arith = "off";

cyclonev_lcell_comb \D_src1_prelim[3]~13 (
	.dataa(!\M_wr_data_unfiltered[3]~8_combout ),
	.datab(!\W_wr_data[3]~q ),
	.datac(!\D_src1_hazard_M~combout ),
	.datad(!\D_src1_hazard_W~combout ),
	.datae(!\processor_cpu_register_bank_a|the_altsyncram|auto_generated|q_b[3] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_prelim[3]~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src1_prelim[3]~13 .extended_lut = "off";
defparam \D_src1_prelim[3]~13 .lut_mask = 64'h7FF7FFFF7FF7FFFF;
defparam \D_src1_prelim[3]~13 .shared_arith = "off";

dffeas \E_src1_prelim[3] (
	.clk(clk_clk),
	.d(\D_src1_prelim[3]~13_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_src1_prelim[3]~q ),
	.prn(vcc));
defparam \E_src1_prelim[3] .is_wysiwyg = "true";
defparam \E_src1_prelim[3] .power_up = "low";

cyclonev_lcell_comb \E_logic_result~12 (
	.dataa(!\E_ctrl_src2_choose_imm~q ),
	.datab(!\E_stb_data[2]~9_combout ),
	.datac(!\E_stb_data[2]~10_combout ),
	.datad(!\E_src2_imm[2]~q ),
	.datae(!\E_src1[2]~24_combout ),
	.dataf(!\E_src1[2]~25_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_logic_result~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_logic_result~12 .extended_lut = "off";
defparam \E_logic_result~12 .lut_mask = 64'h6996966996696996;
defparam \E_logic_result~12 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_prelim[1]~16 (
	.dataa(!\M_wr_data_unfiltered[1]~9_combout ),
	.datab(!\D_src2_hazard_M~combout ),
	.datac(!\D_src2_hazard_W~combout ),
	.datad(!\W_wr_data[1]~q ),
	.datae(!\processor_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[1] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_prelim[1]~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_prelim[1]~16 .extended_lut = "off";
defparam \D_src2_prelim[1]~16 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \D_src2_prelim[1]~16 .shared_arith = "off";

dffeas \E_src2_prelim[1] (
	.clk(clk_clk),
	.d(\D_src2_prelim[1]~16_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_src2_prelim[1]~q ),
	.prn(vcc));
defparam \E_src2_prelim[1] .is_wysiwyg = "true";
defparam \E_src2_prelim[1] .power_up = "low";

cyclonev_lcell_comb \E_arith_src2[1]~12 (
	.dataa(!\E_src2_hazard_M~q ),
	.datab(!\E_ctrl_src2_choose_imm~q ),
	.datac(!\M_wr_data_unfiltered[1]~9_combout ),
	.datad(!\E_src2_prelim[1]~q ),
	.datae(!\E_src2_imm[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_arith_src2[1]~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_arith_src2[1]~12 .extended_lut = "off";
defparam \E_arith_src2[1]~12 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \E_arith_src2[1]~12 .shared_arith = "off";

cyclonev_lcell_comb \E_logic_result~13 (
	.dataa(!\E_stb_data[0]~0_combout ),
	.datab(!\E_stb_data[0]~1_combout ),
	.datac(!\E_ctrl_src2_choose_imm~q ),
	.datad(!\E_src2_imm[0]~q ),
	.datae(!\E_src1[0]~27_combout ),
	.dataf(!\E_src1[0]~28_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_logic_result~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_logic_result~13 .extended_lut = "off";
defparam \E_logic_result~13 .lut_mask = 64'h6996966996696996;
defparam \E_logic_result~13 .shared_arith = "off";

cyclonev_lcell_comb \Add10~130 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_logic_result~13_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\Add10~130_cout ),
	.shareout());
defparam \Add10~130 .extended_lut = "off";
defparam \Add10~130 .lut_mask = 64'h00000000000000FF;
defparam \Add10~130 .shared_arith = "off";

cyclonev_lcell_comb \Add10~126 (
	.dataa(!\E_src1_hazard_M~q ),
	.datab(!\M_wr_data_unfiltered[1]~9_combout ),
	.datac(!\E_arith_src2[1]~12_combout ),
	.datad(!\E_src1_prelim[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add10~130_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\Add10~126_cout ),
	.shareout());
defparam \Add10~126 .extended_lut = "off";
defparam \Add10~126 .lut_mask = 64'h0000000000006996;
defparam \Add10~126 .shared_arith = "off";

cyclonev_lcell_comb \Add10~122 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_logic_result~12_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add10~126_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\Add10~122_cout ),
	.shareout());
defparam \Add10~122 .extended_lut = "off";
defparam \Add10~122 .lut_mask = 64'h00000000000000FF;
defparam \Add10~122 .shared_arith = "off";

cyclonev_lcell_comb \Add10~118 (
	.dataa(!\E_src1_hazard_M~q ),
	.datab(!\M_wr_data_unfiltered[3]~8_combout ),
	.datac(!\E_arith_src2[3]~9_combout ),
	.datad(!\E_src1_prelim[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add10~122_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\Add10~118_cout ),
	.shareout());
defparam \Add10~118 .extended_lut = "off";
defparam \Add10~118 .lut_mask = 64'h0000000000006996;
defparam \Add10~118 .shared_arith = "off";

cyclonev_lcell_comb \Add10~114 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_logic_result~11_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add10~118_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\Add10~114_cout ),
	.shareout());
defparam \Add10~114 .extended_lut = "off";
defparam \Add10~114 .lut_mask = 64'h00000000000000FF;
defparam \Add10~114 .shared_arith = "off";

cyclonev_lcell_comb \Add10~110 (
	.dataa(!\E_src1_hazard_M~q ),
	.datab(!\M_wr_data_unfiltered[5]~0_combout ),
	.datac(!\E_arith_src2[5]~0_combout ),
	.datad(!\E_src1_prelim[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add10~114_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\Add10~110_cout ),
	.shareout());
defparam \Add10~110 .extended_lut = "off";
defparam \Add10~110 .lut_mask = 64'h0000000000006996;
defparam \Add10~110 .shared_arith = "off";

cyclonev_lcell_comb \Add10~106 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_logic_result~10_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add10~110_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\Add10~106_cout ),
	.shareout());
defparam \Add10~106 .extended_lut = "off";
defparam \Add10~106 .lut_mask = 64'h00000000000000FF;
defparam \Add10~106 .shared_arith = "off";

cyclonev_lcell_comb \Add10~102 (
	.dataa(!\E_src1_hazard_M~q ),
	.datab(!\M_wr_data_unfiltered[7]~7_combout ),
	.datac(!\E_arith_src2[7]~8_combout ),
	.datad(!\E_src1_prelim[7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add10~106_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\Add10~102_cout ),
	.shareout());
defparam \Add10~102 .extended_lut = "off";
defparam \Add10~102 .lut_mask = 64'h0000000000006996;
defparam \Add10~102 .shared_arith = "off";

cyclonev_lcell_comb \Add10~98 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_logic_result~9_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add10~102_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\Add10~98_cout ),
	.shareout());
defparam \Add10~98 .extended_lut = "off";
defparam \Add10~98 .lut_mask = 64'h00000000000000FF;
defparam \Add10~98 .shared_arith = "off";

cyclonev_lcell_comb \Add10~94 (
	.dataa(!\E_src1_hazard_M~q ),
	.datab(!\M_wr_data_unfiltered[9]~6_combout ),
	.datac(!\E_arith_src2[9]~7_combout ),
	.datad(!\E_src1_prelim[9]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add10~98_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\Add10~94_cout ),
	.shareout());
defparam \Add10~94 .extended_lut = "off";
defparam \Add10~94 .lut_mask = 64'h0000000000006996;
defparam \Add10~94 .shared_arith = "off";

cyclonev_lcell_comb \Add10~90 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_logic_result~8_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add10~94_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\Add10~90_cout ),
	.shareout());
defparam \Add10~90 .extended_lut = "off";
defparam \Add10~90 .lut_mask = 64'h00000000000000FF;
defparam \Add10~90 .shared_arith = "off";

cyclonev_lcell_comb \Add10~86 (
	.dataa(!\E_src1_hazard_M~q ),
	.datab(!\M_wr_data_unfiltered[11]~5_combout ),
	.datac(!\E_arith_src2[11]~6_combout ),
	.datad(!\E_src1_prelim[11]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add10~90_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\Add10~86_cout ),
	.shareout());
defparam \Add10~86 .extended_lut = "off";
defparam \Add10~86 .lut_mask = 64'h0000000000006996;
defparam \Add10~86 .shared_arith = "off";

cyclonev_lcell_comb \Add10~82 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_logic_result~14_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add10~86_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\Add10~82_cout ),
	.shareout());
defparam \Add10~82 .extended_lut = "off";
defparam \Add10~82 .lut_mask = 64'h00000000000000FF;
defparam \Add10~82 .shared_arith = "off";

cyclonev_lcell_comb \Add10~78 (
	.dataa(!\E_src1_hazard_M~q ),
	.datab(!\M_wr_data_unfiltered[13]~3_combout ),
	.datac(!\E_arith_src2[13]~4_combout ),
	.datad(!\E_src1_prelim[13]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add10~82_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\Add10~78_cout ),
	.shareout());
defparam \Add10~78 .extended_lut = "off";
defparam \Add10~78 .lut_mask = 64'h0000000000006996;
defparam \Add10~78 .shared_arith = "off";

cyclonev_lcell_comb \Add10~74 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_logic_result~18_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add10~78_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\Add10~74_cout ),
	.shareout());
defparam \Add10~74 .extended_lut = "off";
defparam \Add10~74 .lut_mask = 64'h00000000000000FF;
defparam \Add10~74 .shared_arith = "off";

cyclonev_lcell_comb \Add10~70 (
	.dataa(!\E_src1_hazard_M~q ),
	.datab(!\M_wr_data_unfiltered[15]~1_combout ),
	.datac(!\E_arith_src2[15]~2_combout ),
	.datad(!\E_src1_prelim[15]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add10~74_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\Add10~70_cout ),
	.shareout());
defparam \Add10~70 .extended_lut = "off";
defparam \Add10~70 .lut_mask = 64'h0000000000006996;
defparam \Add10~70 .shared_arith = "off";

cyclonev_lcell_comb \Add10~66 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_logic_result~7_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add10~70_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\Add10~66_cout ),
	.shareout());
defparam \Add10~66 .extended_lut = "off";
defparam \Add10~66 .lut_mask = 64'h00000000000000FF;
defparam \Add10~66 .shared_arith = "off";

cyclonev_lcell_comb \Add10~62 (
	.dataa(!\E_src1_hazard_M~q ),
	.datab(!\M_wr_data_unfiltered[17]~18_combout ),
	.datac(!\E_arith_src2[17]~13_combout ),
	.datad(!\E_src1_prelim[17]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add10~66_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\Add10~62_cout ),
	.shareout());
defparam \Add10~62 .extended_lut = "off";
defparam \Add10~62 .lut_mask = 64'h0000000000006996;
defparam \Add10~62 .shared_arith = "off";

cyclonev_lcell_comb \Add10~58 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_logic_result~6_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add10~62_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\Add10~58_cout ),
	.shareout());
defparam \Add10~58 .extended_lut = "off";
defparam \Add10~58 .lut_mask = 64'h00000000000000FF;
defparam \Add10~58 .shared_arith = "off";

cyclonev_lcell_comb \Add10~54 (
	.dataa(!\E_src1_hazard_M~q ),
	.datab(!\M_wr_data_unfiltered[19]~22_combout ),
	.datac(!\E_arith_src2[19]~16_combout ),
	.datad(!\E_src1_prelim[19]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add10~58_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\Add10~54_cout ),
	.shareout());
defparam \Add10~54 .extended_lut = "off";
defparam \Add10~54 .lut_mask = 64'h0000000000006996;
defparam \Add10~54 .shared_arith = "off";

cyclonev_lcell_comb \Add10~50 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_logic_result~5_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add10~54_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\Add10~50_cout ),
	.shareout());
defparam \Add10~50 .extended_lut = "off";
defparam \Add10~50 .lut_mask = 64'h00000000000000FF;
defparam \Add10~50 .shared_arith = "off";

cyclonev_lcell_comb \Add10~46 (
	.dataa(!\E_src1_hazard_M~q ),
	.datab(!\M_wr_data_unfiltered[21]~21_combout ),
	.datac(!\E_arith_src2[21]~15_combout ),
	.datad(!\E_src1_prelim[21]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add10~50_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\Add10~46_cout ),
	.shareout());
defparam \Add10~46 .extended_lut = "off";
defparam \Add10~46 .lut_mask = 64'h0000000000006996;
defparam \Add10~46 .shared_arith = "off";

cyclonev_lcell_comb \Add10~42 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_logic_result~4_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add10~46_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\Add10~42_cout ),
	.shareout());
defparam \Add10~42 .extended_lut = "off";
defparam \Add10~42 .lut_mask = 64'h00000000000000FF;
defparam \Add10~42 .shared_arith = "off";

cyclonev_lcell_comb \Add10~38 (
	.dataa(!\E_src1_hazard_M~q ),
	.datab(!\M_wr_data_unfiltered[23]~24_combout ),
	.datac(!\E_arith_src2[23]~17_combout ),
	.datad(!\E_src1_prelim[23]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add10~42_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\Add10~38_cout ),
	.shareout());
defparam \Add10~38 .extended_lut = "off";
defparam \Add10~38 .lut_mask = 64'h0000000000006996;
defparam \Add10~38 .shared_arith = "off";

cyclonev_lcell_comb \Add10~34 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_logic_result~3_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add10~38_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\Add10~34_cout ),
	.shareout());
defparam \Add10~34 .extended_lut = "off";
defparam \Add10~34 .lut_mask = 64'h00000000000000FF;
defparam \Add10~34 .shared_arith = "off";

cyclonev_lcell_comb \Add10~30 (
	.dataa(!\E_src1_hazard_M~q ),
	.datab(!\M_wr_data_unfiltered[25]~26_combout ),
	.datac(!\E_arith_src2[25]~19_combout ),
	.datad(!\E_src1_prelim[25]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add10~34_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\Add10~30_cout ),
	.shareout());
defparam \Add10~30 .extended_lut = "off";
defparam \Add10~30 .lut_mask = 64'h0000000000006996;
defparam \Add10~30 .shared_arith = "off";

cyclonev_lcell_comb \Add10~26 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_logic_result~2_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add10~30_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\Add10~26_cout ),
	.shareout());
defparam \Add10~26 .extended_lut = "off";
defparam \Add10~26 .lut_mask = 64'h00000000000000FF;
defparam \Add10~26 .shared_arith = "off";

cyclonev_lcell_comb \Add10~22 (
	.dataa(!\E_src1_hazard_M~q ),
	.datab(!\M_wr_data_unfiltered[27]~25_combout ),
	.datac(!\E_arith_src2[27]~18_combout ),
	.datad(!\E_src1_prelim[27]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add10~26_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\Add10~22_cout ),
	.shareout());
defparam \Add10~22 .extended_lut = "off";
defparam \Add10~22 .lut_mask = 64'h0000000000006996;
defparam \Add10~22 .shared_arith = "off";

cyclonev_lcell_comb \Add10~18 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_logic_result~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add10~22_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\Add10~18_cout ),
	.shareout());
defparam \Add10~18 .extended_lut = "off";
defparam \Add10~18 .lut_mask = 64'h00000000000000FF;
defparam \Add10~18 .shared_arith = "off";

cyclonev_lcell_comb \Add10~14 (
	.dataa(!\E_src1_hazard_M~q ),
	.datab(!\M_wr_data_unfiltered[29]~20_combout ),
	.datac(!\E_arith_src2[29]~14_combout ),
	.datad(!\E_src1_prelim[29]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add10~18_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\Add10~14_cout ),
	.shareout());
defparam \Add10~14 .extended_lut = "off";
defparam \Add10~14 .lut_mask = 64'h0000000000006996;
defparam \Add10~14 .shared_arith = "off";

cyclonev_lcell_comb \Add10~10 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_logic_result~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add10~14_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\Add10~10_cout ),
	.shareout());
defparam \Add10~10 .extended_lut = "off";
defparam \Add10~10 .lut_mask = 64'h00000000000000FF;
defparam \Add10~10 .shared_arith = "off";

cyclonev_lcell_comb \Add10~6 (
	.dataa(!\E_src1_hazard_M~q ),
	.datab(!\M_wr_data_unfiltered[31]~17_combout ),
	.datac(!\E_src2[31]~0_combout ),
	.datad(!\E_src1_prelim[31]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add10~10_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\Add10~6_cout ),
	.shareout());
defparam \Add10~6 .extended_lut = "off";
defparam \Add10~6 .lut_mask = 64'h0000000000006996;
defparam \Add10~6 .shared_arith = "off";

cyclonev_lcell_comb \Add10~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add10~6_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add10~1_sumout ),
	.cout(),
	.shareout());
defparam \Add10~1 .extended_lut = "off";
defparam \Add10~1 .lut_mask = 64'h0000000000000000;
defparam \Add10~1 .shared_arith = "off";

cyclonev_lcell_comb \Add8~61 (
	.dataa(gnd),
	.datab(!\E_ctrl_alu_subtract~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add8~74 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add8~61_sumout ),
	.cout(),
	.shareout());
defparam \Add8~61 .extended_lut = "off";
defparam \Add8~61 .lut_mask = 64'h0000000000003333;
defparam \Add8~61 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_break~1 (
	.dataa(!\D_iw[16]~q ),
	.datab(!\D_iw[14]~q ),
	.datac(!\D_ctrl_break~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_break~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_break~1 .extended_lut = "off";
defparam \D_ctrl_break~1 .lut_mask = 64'hDFDFDFDFDFDFDFDF;
defparam \D_ctrl_break~1 .shared_arith = "off";

dffeas E_ctrl_break(
	.clk(clk_clk),
	.d(\D_ctrl_break~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_ctrl_break~q ),
	.prn(vcc));
defparam E_ctrl_break.is_wysiwyg = "true";
defparam E_ctrl_break.power_up = "low";

cyclonev_lcell_comb \D_ctrl_exception~1 (
	.dataa(!\D_iw[11]~q ),
	.datab(!\D_iw[12]~q ),
	.datac(!\D_iw[13]~q ),
	.datad(!\D_iw[14]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_exception~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_exception~1 .extended_lut = "off";
defparam \D_ctrl_exception~1 .lut_mask = 64'hFFDFFFDFFFDFFFDF;
defparam \D_ctrl_exception~1 .shared_arith = "off";

cyclonev_lcell_comb D_ctrl_exception(
	.dataa(!\D_iw[16]~q ),
	.datab(!\D_iw[15]~q ),
	.datac(!\Equal4~0_combout ),
	.datad(!\D_ctrl_exception~1_combout ),
	.datae(!\D_ctrl_exception~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_exception~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam D_ctrl_exception.extended_lut = "off";
defparam D_ctrl_exception.lut_mask = 64'hFFFFDFFFFFFFDFFF;
defparam D_ctrl_exception.shared_arith = "off";

dffeas E_ctrl_exception(
	.clk(clk_clk),
	.d(\D_ctrl_exception~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_ctrl_exception~q ),
	.prn(vcc));
defparam E_ctrl_exception.is_wysiwyg = "true";
defparam E_ctrl_exception.power_up = "low";

cyclonev_lcell_comb \D_ctrl_crst~1 (
	.dataa(!\D_iw[16]~q ),
	.datab(!\D_iw[15]~q ),
	.datac(!\D_iw[14]~q ),
	.datad(!\D_ctrl_crst~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_crst~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_crst~1 .extended_lut = "off";
defparam \D_ctrl_crst~1 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \D_ctrl_crst~1 .shared_arith = "off";

dffeas E_ctrl_crst(
	.clk(clk_clk),
	.d(\D_ctrl_crst~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_ctrl_crst~q ),
	.prn(vcc));
defparam E_ctrl_crst.is_wysiwyg = "true";
defparam E_ctrl_crst.power_up = "low";

dffeas \E_iw[6] (
	.clk(clk_clk),
	.d(\D_iw[6]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_iw[6]~q ),
	.prn(vcc));
defparam \E_iw[6] .is_wysiwyg = "true";
defparam \E_iw[6] .power_up = "low";

dffeas \E_iw[7] (
	.clk(clk_clk),
	.d(\D_iw[7]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_iw[7]~q ),
	.prn(vcc));
defparam \E_iw[7] .is_wysiwyg = "true";
defparam \E_iw[7] .power_up = "low";

dffeas \E_iw[8] (
	.clk(clk_clk),
	.d(\D_iw[8]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_iw[8]~q ),
	.prn(vcc));
defparam \E_iw[8] .is_wysiwyg = "true";
defparam \E_iw[8] .power_up = "low";

cyclonev_lcell_comb \Equal107~2 (
	.dataa(!\D_iw[16]~q ),
	.datab(!\D_iw[15]~q ),
	.datac(!\D_iw[14]~q ),
	.datad(!\D_iw[11]~q ),
	.datae(!\D_ctrl_crst~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal107~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal107~2 .extended_lut = "off";
defparam \Equal107~2 .lut_mask = 64'hFFDFFFFFFFDFFFFF;
defparam \Equal107~2 .shared_arith = "off";

dffeas E_ctrl_wrctl_inst(
	.clk(clk_clk),
	.d(\Equal107~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_ctrl_wrctl_inst~q ),
	.prn(vcc));
defparam E_ctrl_wrctl_inst.is_wysiwyg = "true";
defparam E_ctrl_wrctl_inst.power_up = "low";

cyclonev_lcell_comb \E_op_eret~1 (
	.dataa(!\E_iw[16]~q ),
	.datab(!\E_iw[15]~q ),
	.datac(!\E_iw[13]~q ),
	.datad(!\Equal130~0_combout ),
	.datae(!\E_op_eret~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_op_eret~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_op_eret~1 .extended_lut = "off";
defparam \E_op_eret~1 .lut_mask = 64'hFEFFFFFFFEFFFFFF;
defparam \E_op_eret~1 .shared_arith = "off";

cyclonev_lcell_comb \M_status_reg_pie_inst_nxt~0 (
	.dataa(gnd),
	.datab(!\E_iw[6]~q ),
	.datac(!\E_iw[7]~q ),
	.datad(!\E_iw[8]~q ),
	.datae(!\E_ctrl_wrctl_inst~q ),
	.dataf(!\E_op_eret~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_status_reg_pie_inst_nxt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_status_reg_pie_inst_nxt~0 .extended_lut = "off";
defparam \M_status_reg_pie_inst_nxt~0 .lut_mask = 64'hFFFFFFFFFFFCFFFF;
defparam \M_status_reg_pie_inst_nxt~0 .shared_arith = "off";

cyclonev_lcell_comb E_wrctl_estatus(
	.dataa(!\E_iw[6]~q ),
	.datab(!\E_iw[7]~q ),
	.datac(!\E_iw[8]~q ),
	.datad(!\E_ctrl_wrctl_inst~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_wrctl_estatus~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam E_wrctl_estatus.extended_lut = "off";
defparam E_wrctl_estatus.lut_mask = 64'hFDFFFDFFFDFFFDFF;
defparam E_wrctl_estatus.shared_arith = "off";

cyclonev_lcell_comb \M_estatus_reg_pie_inst_nxt~0 (
	.dataa(!\M_status_reg_pie~q ),
	.datab(!\M_estatus_reg_pie~q ),
	.datac(!\E_ctrl_exception~q ),
	.datad(!\E_ctrl_crst~q ),
	.datae(!\E_wrctl_estatus~combout ),
	.dataf(!\E_wrctl_data_bstatus_reg_pie~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_estatus_reg_pie_inst_nxt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_estatus_reg_pie_inst_nxt~0 .extended_lut = "off";
defparam \M_estatus_reg_pie_inst_nxt~0 .lut_mask = 64'hFF7FFFF7FFFFFFFF;
defparam \M_estatus_reg_pie_inst_nxt~0 .shared_arith = "off";

dffeas M_estatus_reg_pie(
	.clk(clk_clk),
	.d(\M_estatus_reg_pie_inst_nxt~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\M_status_reg_pie~0_combout ),
	.q(\M_estatus_reg_pie~q ),
	.prn(vcc));
defparam M_estatus_reg_pie.is_wysiwyg = "true";
defparam M_estatus_reg_pie.power_up = "low";

cyclonev_lcell_comb E_wrctl_bstatus(
	.dataa(!\E_iw[6]~q ),
	.datab(!\E_iw[7]~q ),
	.datac(!\E_iw[8]~q ),
	.datad(!\E_ctrl_wrctl_inst~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_wrctl_bstatus~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam E_wrctl_bstatus.extended_lut = "off";
defparam E_wrctl_bstatus.lut_mask = 64'hFBFFFBFFFBFFFBFF;
defparam E_wrctl_bstatus.shared_arith = "off";

cyclonev_lcell_comb \M_bstatus_reg_pie_inst_nxt~0 (
	.dataa(!\M_status_reg_pie~q ),
	.datab(!\M_bstatus_reg_pie~q ),
	.datac(!\E_ctrl_break~q ),
	.datad(!\E_wrctl_bstatus~combout ),
	.datae(!\E_wrctl_data_bstatus_reg_pie~2_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_bstatus_reg_pie_inst_nxt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_bstatus_reg_pie_inst_nxt~0 .extended_lut = "off";
defparam \M_bstatus_reg_pie_inst_nxt~0 .lut_mask = 64'h7FF7FFFF7FF7FFFF;
defparam \M_bstatus_reg_pie_inst_nxt~0 .shared_arith = "off";

dffeas M_bstatus_reg_pie(
	.clk(clk_clk),
	.d(\M_bstatus_reg_pie_inst_nxt~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\M_status_reg_pie~0_combout ),
	.q(\M_bstatus_reg_pie~q ),
	.prn(vcc));
defparam M_bstatus_reg_pie.is_wysiwyg = "true";
defparam M_bstatus_reg_pie.power_up = "low";

cyclonev_lcell_comb \M_status_reg_pie_inst_nxt~1 (
	.dataa(!\M_status_reg_pie~q ),
	.datab(!\E_iw[6]~q ),
	.datac(!\E_iw[7]~q ),
	.datad(!\E_iw[8]~q ),
	.datae(!\E_ctrl_wrctl_inst~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_status_reg_pie_inst_nxt~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_status_reg_pie_inst_nxt~1 .extended_lut = "off";
defparam \M_status_reg_pie_inst_nxt~1 .lut_mask = 64'hFFFF7FFFFFFF7FFF;
defparam \M_status_reg_pie_inst_nxt~1 .shared_arith = "off";

cyclonev_lcell_comb \M_status_reg_pie_inst_nxt~2 (
	.dataa(!\E_iw[14]~q ),
	.datab(!\M_estatus_reg_pie~q ),
	.datac(!\M_bstatus_reg_pie~q ),
	.datad(!\E_op_eret~1_combout ),
	.datae(!\M_status_reg_pie_inst_nxt~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_status_reg_pie_inst_nxt~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_status_reg_pie_inst_nxt~2 .extended_lut = "off";
defparam \M_status_reg_pie_inst_nxt~2 .lut_mask = 64'h7FBFFFFF7FBFFFFF;
defparam \M_status_reg_pie_inst_nxt~2 .shared_arith = "off";

cyclonev_lcell_comb \M_status_reg_pie_inst_nxt~3 (
	.dataa(!\E_ctrl_break~q ),
	.datab(!\E_ctrl_exception~q ),
	.datac(!\E_ctrl_crst~q ),
	.datad(!\E_wrctl_data_bstatus_reg_pie~2_combout ),
	.datae(!\M_status_reg_pie_inst_nxt~0_combout ),
	.dataf(!\M_status_reg_pie_inst_nxt~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_status_reg_pie_inst_nxt~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_status_reg_pie_inst_nxt~3 .extended_lut = "off";
defparam \M_status_reg_pie_inst_nxt~3 .lut_mask = 64'hFEFFFFFFFFFFFFFF;
defparam \M_status_reg_pie_inst_nxt~3 .shared_arith = "off";

dffeas M_status_reg_pie(
	.clk(clk_clk),
	.d(\M_status_reg_pie_inst_nxt~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\M_status_reg_pie~0_combout ),
	.q(\M_status_reg_pie~q ),
	.prn(vcc));
defparam M_status_reg_pie.is_wysiwyg = "true";
defparam M_status_reg_pie.power_up = "low";

cyclonev_lcell_comb \D_control_reg_rddata_muxed[0]~1 (
	.dataa(!\D_iw[8]~q ),
	.datab(!\D_iw[7]~q ),
	.datac(!\D_iw[6]~q ),
	.datad(!\M_status_reg_pie~q ),
	.datae(!\M_estatus_reg_pie~q ),
	.dataf(!\M_bstatus_reg_pie~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_control_reg_rddata_muxed[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_control_reg_rddata_muxed[0]~1 .extended_lut = "off";
defparam \D_control_reg_rddata_muxed[0]~1 .lut_mask = 64'hBEFFFFFFFFFFFFFF;
defparam \D_control_reg_rddata_muxed[0]~1 .shared_arith = "off";

dffeas \E_control_reg_rddata[0] (
	.clk(clk_clk),
	.d(\D_control_reg_rddata_muxed[0]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_control_reg_rddata[0]~q ),
	.prn(vcc));
defparam \E_control_reg_rddata[0] .is_wysiwyg = "true";
defparam \E_control_reg_rddata[0] .power_up = "low";

cyclonev_lcell_comb \E_wrctl_data_bstatus_reg_pie~0 (
	.dataa(!\E_ctrl_logic~q ),
	.datab(!\E_src1[0]~29_combout ),
	.datac(!\E_compare_op[1]~q ),
	.datad(!\E_compare_op[0]~q ),
	.datae(!\E_arith_src2[0]~11_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_wrctl_data_bstatus_reg_pie~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_wrctl_data_bstatus_reg_pie~0 .extended_lut = "off";
defparam \E_wrctl_data_bstatus_reg_pie~0 .lut_mask = 64'h7DD7D77D7DD7D77D;
defparam \E_wrctl_data_bstatus_reg_pie~0 .shared_arith = "off";

cyclonev_lcell_comb \E_wrctl_data_bstatus_reg_pie~1 (
	.dataa(!\E_ctrl_rdctl_inst~q ),
	.datab(!\E_alu_result~0_combout ),
	.datac(!\E_control_reg_rddata[0]~q ),
	.datad(!\Add8~65_sumout ),
	.datae(!\E_wrctl_data_bstatus_reg_pie~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_wrctl_data_bstatus_reg_pie~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_wrctl_data_bstatus_reg_pie~1 .extended_lut = "off";
defparam \E_wrctl_data_bstatus_reg_pie~1 .lut_mask = 64'hFFFFFFFEFFFFFFFE;
defparam \E_wrctl_data_bstatus_reg_pie~1 .shared_arith = "off";

cyclonev_lcell_comb \E_wrctl_data_bstatus_reg_pie~2 (
	.dataa(!\E_ctrl_cmp~q ),
	.datab(!\E_compare_op[1]~q ),
	.datac(!\E_compare_op[0]~q ),
	.datad(!\Add10~1_sumout ),
	.datae(!\Add8~61_sumout ),
	.dataf(!\E_wrctl_data_bstatus_reg_pie~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_wrctl_data_bstatus_reg_pie~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_wrctl_data_bstatus_reg_pie~2 .extended_lut = "off";
defparam \E_wrctl_data_bstatus_reg_pie~2 .lut_mask = 64'hFFFFFFFF7DD7D77D;
defparam \E_wrctl_data_bstatus_reg_pie~2 .shared_arith = "off";

dffeas \M_alu_result[0] (
	.clk(clk_clk),
	.d(\E_wrctl_data_bstatus_reg_pie~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\M_alu_result[0]~q ),
	.prn(vcc));
defparam \M_alu_result[0] .is_wysiwyg = "true";
defparam \M_alu_result[0] .power_up = "low";

cyclonev_lcell_comb M_ld_align_sh8(
	.dataa(!\M_alu_result[0]~q ),
	.datab(!\Equal2~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_ld_align_sh8~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam M_ld_align_sh8.extended_lut = "off";
defparam M_ld_align_sh8.lut_mask = 64'h7777777777777777;
defparam M_ld_align_sh8.shared_arith = "off";

cyclonev_lcell_comb \av_ld_byte0_data[1]~7 (
	.dataa(!\d_readdata_d1[1]~q ),
	.datab(!\d_readdata_d1[17]~q ),
	.datac(!\d_readdata_d1[9]~q ),
	.datad(!\d_readdata_d1[25]~q ),
	.datae(!\M_ld_align_sh16~combout ),
	.dataf(!\M_ld_align_sh8~combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_ld_byte0_data[1]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_ld_byte0_data[1]~7 .extended_lut = "off";
defparam \av_ld_byte0_data[1]~7 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \av_ld_byte0_data[1]~7 .shared_arith = "off";

dffeas \av_ld_data_aligned_or_div[1] (
	.clk(clk_clk),
	.d(\av_ld_byte0_data[1]~7_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\av_ld_data_aligned_or_div[1]~q ),
	.prn(vcc));
defparam \av_ld_data_aligned_or_div[1] .is_wysiwyg = "true";
defparam \av_ld_data_aligned_or_div[1] .power_up = "low";

cyclonev_lcell_comb \M_wr_data_unfiltered[1]~9 (
	.dataa(!\M_ctrl_shift_rot~q ),
	.datab(!\av_ld_or_div_done~q ),
	.datac(!\M_shift_rot_result[1]~q ),
	.datad(!\av_ld_data_aligned_or_div[1]~q ),
	.datae(!\M_alu_result[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_wr_data_unfiltered[1]~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_wr_data_unfiltered[1]~9 .extended_lut = "off";
defparam \M_wr_data_unfiltered[1]~9 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \M_wr_data_unfiltered[1]~9 .shared_arith = "off";

cyclonev_lcell_comb \E_stb_data[1]~12 (
	.dataa(!\E_src2_hazard_M~q ),
	.datab(!\M_wr_data_unfiltered[1]~9_combout ),
	.datac(!\E_src2_prelim[1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_stb_data[1]~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_stb_data[1]~12 .extended_lut = "off";
defparam \E_stb_data[1]~12 .lut_mask = 64'h2727272727272727;
defparam \E_stb_data[1]~12 .shared_arith = "off";

cyclonev_lcell_comb \M_ienable_reg_irq16~1 (
	.dataa(!\E_iw[6]~q ),
	.datab(!\E_iw[7]~q ),
	.datac(!\E_iw[8]~q ),
	.datad(!\E_ctrl_wrctl_inst~q ),
	.datae(!\W_stall~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_ienable_reg_irq16~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_ienable_reg_irq16~1 .extended_lut = "off";
defparam \M_ienable_reg_irq16~1 .lut_mask = 64'hF7FFFFFFF7FFFFFF;
defparam \M_ienable_reg_irq16~1 .shared_arith = "off";

cyclonev_lcell_comb \M_ienable_reg_irq16~0 (
	.dataa(!d_write1),
	.datab(!d_read1),
	.datac(!WideOr1),
	.datad(!read_accepted),
	.datae(!\E_valid~1_combout ),
	.dataf(!\M_ienable_reg_irq16~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_ienable_reg_irq16~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_ienable_reg_irq16~0 .extended_lut = "off";
defparam \M_ienable_reg_irq16~0 .lut_mask = 64'hB8FFFFFFFFFFFFFF;
defparam \M_ienable_reg_irq16~0 .shared_arith = "off";

dffeas M_ienable_reg_irq1(
	.clk(clk_clk),
	.d(\E_wrctl_data_ienable_reg_irq1~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\M_ienable_reg_irq16~0_combout ),
	.q(\M_ienable_reg_irq1~q ),
	.prn(vcc));
defparam M_ienable_reg_irq1.is_wysiwyg = "true";
defparam M_ienable_reg_irq1.power_up = "low";

cyclonev_lcell_comb M_ipending_reg_irq1_nxt(
	.dataa(!\M_ienable_reg_irq1~q ),
	.datab(!\the_processor_cpu_nios2_oci|the_processor_cpu_nios2_avalon_reg|oci_ienable[1]~q ),
	.datac(!timeout_occurred),
	.datad(!control_register_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_ipending_reg_irq1_nxt~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam M_ipending_reg_irq1_nxt.extended_lut = "off";
defparam M_ipending_reg_irq1_nxt.lut_mask = 64'hDFFFDFFFDFFFDFFF;
defparam M_ipending_reg_irq1_nxt.shared_arith = "off";

dffeas M_ipending_reg_irq1(
	.clk(clk_clk),
	.d(\M_ipending_reg_irq1_nxt~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\M_ipending_reg_irq1~q ),
	.prn(vcc));
defparam M_ipending_reg_irq1.is_wysiwyg = "true";
defparam M_ipending_reg_irq1.power_up = "low";

cyclonev_lcell_comb \D_control_reg_rddata_muxed[1]~2 (
	.dataa(!\D_iw[8]~q ),
	.datab(!\D_iw[7]~q ),
	.datac(!\D_iw[6]~q ),
	.datad(!\M_ipending_reg_irq1~q ),
	.datae(!\M_ienable_reg_irq1~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_control_reg_rddata_muxed[1]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_control_reg_rddata_muxed[1]~2 .extended_lut = "off";
defparam \D_control_reg_rddata_muxed[1]~2 .lut_mask = 64'h96FFFFFF96FFFFFF;
defparam \D_control_reg_rddata_muxed[1]~2 .shared_arith = "off";

dffeas \E_control_reg_rddata[1] (
	.clk(clk_clk),
	.d(\D_control_reg_rddata_muxed[1]~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_control_reg_rddata[1]~q ),
	.prn(vcc));
defparam \E_control_reg_rddata[1] .is_wysiwyg = "true";
defparam \E_control_reg_rddata[1] .power_up = "low";

cyclonev_lcell_comb \E_wrctl_data_ienable_reg_irq1~0 (
	.dataa(!\E_ctrl_logic~q ),
	.datab(!\E_src1[1]~30_combout ),
	.datac(!\E_compare_op[1]~q ),
	.datad(!\E_compare_op[0]~q ),
	.datae(!\E_arith_src2[1]~12_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_wrctl_data_ienable_reg_irq1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_wrctl_data_ienable_reg_irq1~0 .extended_lut = "off";
defparam \E_wrctl_data_ienable_reg_irq1~0 .lut_mask = 64'h7DD7D77D7DD7D77D;
defparam \E_wrctl_data_ienable_reg_irq1~0 .shared_arith = "off";

cyclonev_lcell_comb \E_wrctl_data_ienable_reg_irq1~1 (
	.dataa(!\E_ctrl_rdctl_inst~q ),
	.datab(!\E_alu_result~0_combout ),
	.datac(!\Add8~69_sumout ),
	.datad(!\E_control_reg_rddata[1]~q ),
	.datae(!\E_wrctl_data_ienable_reg_irq1~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_wrctl_data_ienable_reg_irq1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_wrctl_data_ienable_reg_irq1~1 .extended_lut = "off";
defparam \E_wrctl_data_ienable_reg_irq1~1 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \E_wrctl_data_ienable_reg_irq1~1 .shared_arith = "off";

dffeas \M_alu_result[1] (
	.clk(clk_clk),
	.d(\E_wrctl_data_ienable_reg_irq1~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\M_alu_result[1]~q ),
	.prn(vcc));
defparam \M_alu_result[1] .is_wysiwyg = "true";
defparam \M_alu_result[1] .power_up = "low";

cyclonev_lcell_comb M_ld_align_sh16(
	.dataa(!\M_alu_result[1]~q ),
	.datab(!\M_iw[4]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_ld_align_sh16~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam M_ld_align_sh16.extended_lut = "off";
defparam M_ld_align_sh16.lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam M_ld_align_sh16.shared_arith = "off";

cyclonev_lcell_comb \av_ld_byte0_data[3]~5 (
	.dataa(!\d_readdata_d1[3]~q ),
	.datab(!\d_readdata_d1[19]~q ),
	.datac(!\d_readdata_d1[11]~q ),
	.datad(!\d_readdata_d1[27]~q ),
	.datae(!\M_ld_align_sh16~combout ),
	.dataf(!\M_ld_align_sh8~combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_ld_byte0_data[3]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_ld_byte0_data[3]~5 .extended_lut = "off";
defparam \av_ld_byte0_data[3]~5 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \av_ld_byte0_data[3]~5 .shared_arith = "off";

dffeas \av_ld_data_aligned_or_div[3] (
	.clk(clk_clk),
	.d(\av_ld_byte0_data[3]~5_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\av_ld_data_aligned_or_div[3]~q ),
	.prn(vcc));
defparam \av_ld_data_aligned_or_div[3] .is_wysiwyg = "true";
defparam \av_ld_data_aligned_or_div[3] .power_up = "low";

cyclonev_lcell_comb \M_wr_data_unfiltered[3]~8 (
	.dataa(!M_alu_result_3),
	.datab(!\M_ctrl_shift_rot~q ),
	.datac(!\av_ld_or_div_done~q ),
	.datad(!\M_shift_rot_result[3]~q ),
	.datae(!\av_ld_data_aligned_or_div[3]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_wr_data_unfiltered[3]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_wr_data_unfiltered[3]~8 .extended_lut = "off";
defparam \M_wr_data_unfiltered[3]~8 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \M_wr_data_unfiltered[3]~8 .shared_arith = "off";

cyclonev_lcell_comb \E_src1[3]~23 (
	.dataa(!\M_wr_data_unfiltered[3]~8_combout ),
	.datab(!\E_src1_hazard_M~q ),
	.datac(!\E_src1_prelim[3]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_src1[3]~23_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_src1[3]~23 .extended_lut = "off";
defparam \E_src1[3]~23 .lut_mask = 64'h4747474747474747;
defparam \E_src1[3]~23 .shared_arith = "off";

cyclonev_lcell_comb \M_shift_rot_result_nxt[3]~14 (
	.dataa(!\M_shift_rot_stall~q ),
	.datab(!\E_src1[3]~23_combout ),
	.datac(!\M_shift_rot_result[2]~q ),
	.datad(!\M_shift_rot_result[4]~q ),
	.datae(!\M_ctrl_shift_rot_right~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_shift_rot_result_nxt[3]~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_shift_rot_result_nxt[3]~14 .extended_lut = "off";
defparam \M_shift_rot_result_nxt[3]~14 .lut_mask = 64'h7FFFBFFF7FFFBFFF;
defparam \M_shift_rot_result_nxt[3]~14 .shared_arith = "off";

dffeas \M_shift_rot_result[3] (
	.clk(clk_clk),
	.d(\M_shift_rot_result_nxt[3]~14_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\M_shift_rot_result[3]~q ),
	.prn(vcc));
defparam \M_shift_rot_result[3] .is_wysiwyg = "true";
defparam \M_shift_rot_result[3] .power_up = "low";

cyclonev_lcell_comb \M_shift_rot_result_nxt[2]~15 (
	.dataa(!\M_shift_rot_stall~q ),
	.datab(!\M_shift_rot_result[3]~q ),
	.datac(!\E_src1[2]~26_combout ),
	.datad(!\M_shift_rot_result[1]~q ),
	.datae(!\M_ctrl_shift_rot_right~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_shift_rot_result_nxt[2]~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_shift_rot_result_nxt[2]~15 .extended_lut = "off";
defparam \M_shift_rot_result_nxt[2]~15 .lut_mask = 64'h7FFFBFFF7FFFBFFF;
defparam \M_shift_rot_result_nxt[2]~15 .shared_arith = "off";

dffeas \M_shift_rot_result[2] (
	.clk(clk_clk),
	.d(\M_shift_rot_result_nxt[2]~15_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\M_shift_rot_result[2]~q ),
	.prn(vcc));
defparam \M_shift_rot_result[2] .is_wysiwyg = "true";
defparam \M_shift_rot_result[2] .power_up = "low";

cyclonev_lcell_comb \M_shift_rot_result_nxt[1]~16 (
	.dataa(!\M_shift_rot_result[0]~q ),
	.datab(!\M_shift_rot_stall~q ),
	.datac(!\M_shift_rot_result[2]~q ),
	.datad(!\E_src1[1]~30_combout ),
	.datae(!\M_ctrl_shift_rot_right~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_shift_rot_result_nxt[1]~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_shift_rot_result_nxt[1]~16 .extended_lut = "off";
defparam \M_shift_rot_result_nxt[1]~16 .lut_mask = 64'h7FFFDFFF7FFFDFFF;
defparam \M_shift_rot_result_nxt[1]~16 .shared_arith = "off";

dffeas \M_shift_rot_result[1] (
	.clk(clk_clk),
	.d(\M_shift_rot_result_nxt[1]~16_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\M_shift_rot_result[1]~q ),
	.prn(vcc));
defparam \M_shift_rot_result[1] .is_wysiwyg = "true";
defparam \M_shift_rot_result[1] .power_up = "low";

cyclonev_lcell_comb \M_shift_rot_result_nxt[0]~0 (
	.dataa(!\M_shift_rot_stall~q ),
	.datab(!\M_shift_rot_result[1]~q ),
	.datac(!\E_src1[0]~29_combout ),
	.datad(!\M_ctrl_shift_rot_right~q ),
	.datae(!\M_shift_rot_fill_bit~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_shift_rot_result_nxt[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_shift_rot_result_nxt[0]~0 .extended_lut = "off";
defparam \M_shift_rot_result_nxt[0]~0 .lut_mask = 64'h7FBFFFFF7FBFFFFF;
defparam \M_shift_rot_result_nxt[0]~0 .shared_arith = "off";

dffeas \M_shift_rot_result[0] (
	.clk(clk_clk),
	.d(\M_shift_rot_result_nxt[0]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\M_shift_rot_result[0]~q ),
	.prn(vcc));
defparam \M_shift_rot_result[0] .is_wysiwyg = "true";
defparam \M_shift_rot_result[0] .power_up = "low";

cyclonev_lcell_comb \M_wr_data_unfiltered[0]~10 (
	.dataa(!\M_shift_rot_result[0]~q ),
	.datab(!\M_ctrl_shift_rot~q ),
	.datac(!\av_ld_data_aligned_or_div[0]~q ),
	.datad(!\av_ld_or_div_done~q ),
	.datae(!\M_alu_result[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_wr_data_unfiltered[0]~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_wr_data_unfiltered[0]~10 .extended_lut = "off";
defparam \M_wr_data_unfiltered[0]~10 .lut_mask = 64'h7FDFFFFF7FDFFFFF;
defparam \M_wr_data_unfiltered[0]~10 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_prelim[0]~0 (
	.dataa(!\M_wr_data_unfiltered[0]~10_combout ),
	.datab(!\D_src2_hazard_M~combout ),
	.datac(!\W_wr_data[0]~q ),
	.datad(!\D_src2_hazard_W~combout ),
	.datae(!\processor_cpu_register_bank_b|the_altsyncram|auto_generated|q_b[0] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_prelim[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_prelim[0]~0 .extended_lut = "off";
defparam \D_src2_prelim[0]~0 .lut_mask = 64'h7FDFFFFF7FDFFFFF;
defparam \D_src2_prelim[0]~0 .shared_arith = "off";

dffeas \E_src2_prelim[0] (
	.clk(clk_clk),
	.d(\D_src2_prelim[0]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_src2_prelim[0]~q ),
	.prn(vcc));
defparam \E_src2_prelim[0] .is_wysiwyg = "true";
defparam \E_src2_prelim[0] .power_up = "low";

cyclonev_lcell_comb \E_stb_data[0]~1 (
	.dataa(!\E_src2_hazard_M~q ),
	.datab(!\E_src2_prelim[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_stb_data[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_stb_data[0]~1 .extended_lut = "off";
defparam \E_stb_data[0]~1 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \E_stb_data[0]~1 .shared_arith = "off";

cyclonev_lcell_comb \E_arith_src2[0]~11 (
	.dataa(!\E_ctrl_src2_choose_imm~q ),
	.datab(!\E_src2_imm[0]~q ),
	.datac(!\E_stb_data[0]~0_combout ),
	.datad(!\E_stb_data[0]~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_arith_src2[0]~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_arith_src2[0]~11 .extended_lut = "off";
defparam \E_arith_src2[0]~11 .lut_mask = 64'hFFD8FFD8FFD8FFD8;
defparam \E_arith_src2[0]~11 .shared_arith = "off";

dffeas \M_shift_rot_cnt[0] (
	.clk(clk_clk),
	.d(\M_shift_rot_cnt_nxt[0]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\M_shift_rot_cnt[0]~q ),
	.prn(vcc));
defparam \M_shift_rot_cnt[0] .is_wysiwyg = "true";
defparam \M_shift_rot_cnt[0] .power_up = "low";

cyclonev_lcell_comb \M_shift_rot_cnt_nxt[0]~0 (
	.dataa(!\M_shift_rot_stall~q ),
	.datab(!\E_arith_src2[0]~11_combout ),
	.datac(!\M_shift_rot_cnt[0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_shift_rot_cnt_nxt[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_shift_rot_cnt_nxt[0]~0 .extended_lut = "off";
defparam \M_shift_rot_cnt_nxt[0]~0 .lut_mask = 64'hD8D8D8D8D8D8D8D8;
defparam \M_shift_rot_cnt_nxt[0]~0 .shared_arith = "off";

dffeas \M_shift_rot_cnt[1] (
	.clk(clk_clk),
	.d(\M_shift_rot_cnt_nxt[1]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\M_shift_rot_cnt[1]~q ),
	.prn(vcc));
defparam \M_shift_rot_cnt[1] .is_wysiwyg = "true";
defparam \M_shift_rot_cnt[1] .power_up = "low";

cyclonev_lcell_comb \M_shift_rot_cnt_nxt[1]~1 (
	.dataa(!\M_shift_rot_stall~q ),
	.datab(!\E_arith_src2[1]~12_combout ),
	.datac(!\M_shift_rot_cnt[1]~q ),
	.datad(!\M_shift_rot_cnt[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_shift_rot_cnt_nxt[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_shift_rot_cnt_nxt[1]~1 .extended_lut = "off";
defparam \M_shift_rot_cnt_nxt[1]~1 .lut_mask = 64'hB77BB77BB77BB77B;
defparam \M_shift_rot_cnt_nxt[1]~1 .shared_arith = "off";

cyclonev_lcell_comb \E_arith_src2[2]~10 (
	.dataa(!\E_ctrl_src2_choose_imm~q ),
	.datab(!\E_stb_data[2]~11_combout ),
	.datac(!\E_src2_imm[2]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_arith_src2[2]~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_arith_src2[2]~10 .extended_lut = "off";
defparam \E_arith_src2[2]~10 .lut_mask = 64'h2727272727272727;
defparam \E_arith_src2[2]~10 .shared_arith = "off";

dffeas \M_shift_rot_cnt[2] (
	.clk(clk_clk),
	.d(\M_shift_rot_cnt_nxt[2]~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\M_shift_rot_cnt[2]~q ),
	.prn(vcc));
defparam \M_shift_rot_cnt[2] .is_wysiwyg = "true";
defparam \M_shift_rot_cnt[2] .power_up = "low";

cyclonev_lcell_comb \M_shift_rot_cnt_nxt[2]~2 (
	.dataa(!\M_shift_rot_stall~q ),
	.datab(!\E_arith_src2[2]~10_combout ),
	.datac(!\M_shift_rot_cnt[1]~q ),
	.datad(!\M_shift_rot_cnt[0]~q ),
	.datae(!\M_shift_rot_cnt[2]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_shift_rot_cnt_nxt[2]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_shift_rot_cnt_nxt[2]~2 .extended_lut = "off";
defparam \M_shift_rot_cnt_nxt[2]~2 .lut_mask = 64'h7BB7B77B7BB7B77B;
defparam \M_shift_rot_cnt_nxt[2]~2 .shared_arith = "off";

cyclonev_lcell_comb \E_arith_src2[4]~1 (
	.dataa(!\E_ctrl_src2_choose_imm~q ),
	.datab(!\E_stb_data[4]~5_combout ),
	.datac(!\E_src2_imm[4]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_arith_src2[4]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_arith_src2[4]~1 .extended_lut = "off";
defparam \E_arith_src2[4]~1 .lut_mask = 64'h2727272727272727;
defparam \E_arith_src2[4]~1 .shared_arith = "off";

dffeas \M_shift_rot_cnt[4] (
	.clk(clk_clk),
	.d(\M_shift_rot_cnt_nxt[4]~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\M_shift_rot_cnt[4]~q ),
	.prn(vcc));
defparam \M_shift_rot_cnt[4] .is_wysiwyg = "true";
defparam \M_shift_rot_cnt[4] .power_up = "low";

cyclonev_lcell_comb \Add9~0 (
	.dataa(!\M_shift_rot_cnt[1]~q ),
	.datab(!\M_shift_rot_cnt[0]~q ),
	.datac(!\M_shift_rot_cnt[2]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add9~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add9~0 .extended_lut = "off";
defparam \Add9~0 .lut_mask = 64'hFEFEFEFEFEFEFEFE;
defparam \Add9~0 .shared_arith = "off";

cyclonev_lcell_comb \M_shift_rot_cnt_nxt[3]~4 (
	.dataa(!\M_shift_rot_stall~q ),
	.datab(!\E_arith_src2[3]~9_combout ),
	.datac(!\M_shift_rot_cnt[3]~q ),
	.datad(!\Add9~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_shift_rot_cnt_nxt[3]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_shift_rot_cnt_nxt[3]~4 .extended_lut = "off";
defparam \M_shift_rot_cnt_nxt[3]~4 .lut_mask = 64'hB77BB77BB77BB77B;
defparam \M_shift_rot_cnt_nxt[3]~4 .shared_arith = "off";

dffeas \M_shift_rot_cnt[3] (
	.clk(clk_clk),
	.d(\M_shift_rot_cnt_nxt[3]~4_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\M_shift_rot_cnt[3]~q ),
	.prn(vcc));
defparam \M_shift_rot_cnt[3] .is_wysiwyg = "true";
defparam \M_shift_rot_cnt[3] .power_up = "low";

cyclonev_lcell_comb \M_shift_rot_cnt_nxt[4]~3 (
	.dataa(!\M_shift_rot_stall~q ),
	.datab(!\E_arith_src2[4]~1_combout ),
	.datac(!\M_shift_rot_cnt[4]~q ),
	.datad(!\M_shift_rot_cnt[3]~q ),
	.datae(!\Add9~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_shift_rot_cnt_nxt[4]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_shift_rot_cnt_nxt[4]~3 .extended_lut = "off";
defparam \M_shift_rot_cnt_nxt[4]~3 .lut_mask = 64'h7BB7B77B7BB7B77B;
defparam \M_shift_rot_cnt_nxt[4]~3 .shared_arith = "off";

cyclonev_lcell_comb \Equal198~0 (
	.dataa(!\M_shift_rot_cnt_nxt[1]~1_combout ),
	.datab(!\M_shift_rot_cnt_nxt[2]~2_combout ),
	.datac(!\M_shift_rot_cnt_nxt[4]~3_combout ),
	.datad(!\M_shift_rot_cnt_nxt[3]~4_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal198~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal198~0 .extended_lut = "off";
defparam \Equal198~0 .lut_mask = 64'hFFFEFFFEFFFEFFFE;
defparam \Equal198~0 .shared_arith = "off";

cyclonev_lcell_comb \M_shift_rot_stall_nxt~0 (
	.dataa(!\M_shift_rot_stall~q ),
	.datab(!\M_status_reg_pie~0_combout ),
	.datac(!\E_ctrl_shift_rot~q ),
	.datad(!\M_shift_rot_cnt_nxt[0]~0_combout ),
	.datae(!\Equal198~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_shift_rot_stall_nxt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_shift_rot_stall_nxt~0 .extended_lut = "off";
defparam \M_shift_rot_stall_nxt~0 .lut_mask = 64'hFFFF7FFFFFFF7FFF;
defparam \M_shift_rot_stall_nxt~0 .shared_arith = "off";

dffeas M_shift_rot_stall(
	.clk(clk_clk),
	.d(\M_shift_rot_stall_nxt~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\M_shift_rot_stall~q ),
	.prn(vcc));
defparam M_shift_rot_stall.is_wysiwyg = "true";
defparam M_shift_rot_stall.power_up = "low";

cyclonev_lcell_comb \W_stall~0 (
	.dataa(!\av_ld_or_div_done~q ),
	.datab(!\M_valid_from_E~q ),
	.datac(!\M_ctrl_ld~q ),
	.datad(!\M_shift_rot_stall~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\W_stall~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \W_stall~0 .extended_lut = "off";
defparam \W_stall~0 .lut_mask = 64'hFFFDFFFDFFFDFFFD;
defparam \W_stall~0 .shared_arith = "off";

cyclonev_lcell_comb W_stall(
	.dataa(!d_write1),
	.datab(!d_read1),
	.datac(!WideOr1),
	.datad(!read_accepted),
	.datae(!\W_stall~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\W_stall~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam W_stall.extended_lut = "off";
defparam W_stall.lut_mask = 64'hB8FFFFFFB8FFFFFF;
defparam W_stall.shared_arith = "off";

dffeas \D_iw[14] (
	.clk(clk_clk),
	.d(\F_iw[14]~12_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\F_iw~1_combout ),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\D_iw[14]~q ),
	.prn(vcc));
defparam \D_iw[14] .is_wysiwyg = "true";
defparam \D_iw[14] .power_up = "low";

dffeas \E_iw[14] (
	.clk(clk_clk),
	.d(\D_iw[14]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_iw[14]~q ),
	.prn(vcc));
defparam \E_iw[14] .is_wysiwyg = "true";
defparam \E_iw[14] .power_up = "low";

cyclonev_lcell_comb E_hbreak_req(
	.dataa(!\E_iw[14]~q ),
	.datab(!\E_valid~0_combout ),
	.datac(!\Equal130~0_combout ),
	.datad(!\E_op_eret~0_combout ),
	.datae(!\E_hbreak_req~0_combout ),
	.dataf(!\hbreak_req~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_hbreak_req~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam E_hbreak_req.extended_lut = "off";
defparam E_hbreak_req.lut_mask = 64'hFFFFFFFDFFFFFFFF;
defparam E_hbreak_req.shared_arith = "off";

dffeas \E_iw[21] (
	.clk(clk_clk),
	.d(\D_iw[21]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_iw[21]~q ),
	.prn(vcc));
defparam \E_iw[21] .is_wysiwyg = "true";
defparam \E_iw[21] .power_up = "low";

cyclonev_lcell_comb \E_br_mispredict~0 (
	.dataa(!\E_compare_op[1]~q ),
	.datab(!\E_compare_op[0]~q ),
	.datac(!\Add10~1_sumout ),
	.datad(!\Add8~61_sumout ),
	.datae(!\E_iw[21]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_br_mispredict~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_br_mispredict~0 .extended_lut = "off";
defparam \E_br_mispredict~0 .lut_mask = 64'h9669699696696996;
defparam \E_br_mispredict~0 .shared_arith = "off";

cyclonev_lcell_comb \E_ctrl_br_cond_nxt~0 (
	.dataa(!\D_iw[4]~q ),
	.datab(!\D_iw[5]~q ),
	.datac(!\D_iw[2]~q ),
	.datad(!\D_iw[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_ctrl_br_cond_nxt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_ctrl_br_cond_nxt~0 .extended_lut = "off";
defparam \E_ctrl_br_cond_nxt~0 .lut_mask = 64'hFFD8FFD8FFD8FFD8;
defparam \E_ctrl_br_cond_nxt~0 .shared_arith = "off";

cyclonev_lcell_comb \E_ctrl_br_cond_nxt~1 (
	.dataa(!\D_iw[0]~q ),
	.datab(!\D_iw[1]~q ),
	.datac(!\E_ctrl_br_cond_nxt~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_ctrl_br_cond_nxt~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_ctrl_br_cond_nxt~1 .extended_lut = "off";
defparam \E_ctrl_br_cond_nxt~1 .lut_mask = 64'hFBFBFBFBFBFBFBFB;
defparam \E_ctrl_br_cond_nxt~1 .shared_arith = "off";

dffeas E_ctrl_br_cond(
	.clk(clk_clk),
	.d(\E_ctrl_br_cond_nxt~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_ctrl_br_cond~q ),
	.prn(vcc));
defparam E_ctrl_br_cond.is_wysiwyg = "true";
defparam E_ctrl_br_cond.power_up = "low";

cyclonev_lcell_comb \Equal4~11 (
	.dataa(!\D_iw[0]~q ),
	.datab(!\D_iw[1]~q ),
	.datac(!\D_iw[2]~q ),
	.datad(!\D_iw[3]~q ),
	.datae(!\D_iw[4]~q ),
	.dataf(!\D_iw[5]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal4~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal4~11 .extended_lut = "off";
defparam \Equal4~11 .lut_mask = 64'hFFFFFFFFFFFFFFFD;
defparam \Equal4~11 .shared_arith = "off";

cyclonev_lcell_comb \Equal4~13 (
	.dataa(!\D_iw[0]~q ),
	.datab(!\D_iw[1]~q ),
	.datac(!\D_iw[2]~q ),
	.datad(!\D_iw[3]~q ),
	.datae(!\D_iw[4]~q ),
	.dataf(!\D_iw[5]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal4~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal4~13 .extended_lut = "off";
defparam \Equal4~13 .lut_mask = 64'hFFFFFFFFFFFFFFFE;
defparam \Equal4~13 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_flush_pipe_always~1 (
	.dataa(!\D_iw[14]~q ),
	.datab(!\D_iw[13]~q ),
	.datac(!\D_iw[16]~q ),
	.datad(!\D_iw[11]~q ),
	.datae(!\D_iw[15]~q ),
	.dataf(!\D_iw[12]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_flush_pipe_always~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_flush_pipe_always~1 .extended_lut = "off";
defparam \D_ctrl_flush_pipe_always~1 .lut_mask = 64'hB77B7BB77BB7B77B;
defparam \D_ctrl_flush_pipe_always~1 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_flush_pipe_always~0 (
	.dataa(!\Equal4~0_combout ),
	.datab(!\Equal4~11_combout ),
	.datac(!\Equal4~13_combout ),
	.datad(!\D_ctrl_flush_pipe_always~1_combout ),
	.datae(!\D_ctrl_exception~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_flush_pipe_always~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_flush_pipe_always~0 .extended_lut = "off";
defparam \D_ctrl_flush_pipe_always~0 .lut_mask = 64'hFFFF7FFFFFFF7FFF;
defparam \D_ctrl_flush_pipe_always~0 .shared_arith = "off";

dffeas E_ctrl_flush_pipe_always(
	.clk(clk_clk),
	.d(\D_ctrl_flush_pipe_always~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_ctrl_flush_pipe_always~q ),
	.prn(vcc));
defparam E_ctrl_flush_pipe_always.is_wysiwyg = "true";
defparam E_ctrl_flush_pipe_always.power_up = "low";

cyclonev_lcell_comb \M_pipe_flush_nxt~0 (
	.dataa(!\E_valid~0_combout ),
	.datab(!\E_hbreak_req~combout ),
	.datac(!\E_br_mispredict~0_combout ),
	.datad(!\E_ctrl_br_cond~q ),
	.datae(!\E_ctrl_flush_pipe_always~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_pipe_flush_nxt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_pipe_flush_nxt~0 .extended_lut = "off";
defparam \M_pipe_flush_nxt~0 .lut_mask = 64'hFFFFFFFEFFFFFFFE;
defparam \M_pipe_flush_nxt~0 .shared_arith = "off";

dffeas M_pipe_flush(
	.clk(clk_clk),
	.d(\M_pipe_flush_nxt~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\M_pipe_flush~q ),
	.prn(vcc));
defparam M_pipe_flush.is_wysiwyg = "true";
defparam M_pipe_flush.power_up = "low";

cyclonev_lcell_comb \D_ctrl_br~0 (
	.dataa(!\D_iw[0]~q ),
	.datab(!\D_iw[1]~q ),
	.datac(!\D_iw[2]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_br~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_br~0 .extended_lut = "off";
defparam \D_ctrl_br~0 .lut_mask = 64'hBFBFBFBFBFBFBFBF;
defparam \D_ctrl_br~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal4~12 (
	.dataa(!\D_iw[0]~q ),
	.datab(!\D_iw[1]~q ),
	.datac(!\D_iw[2]~q ),
	.datad(!\D_iw[3]~q ),
	.datae(!\D_iw[4]~q ),
	.dataf(!\D_iw[5]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal4~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal4~12 .extended_lut = "off";
defparam \Equal4~12 .lut_mask = 64'hFFFFFFFFFFFFFFBF;
defparam \Equal4~12 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_jmp_indirect~0 (
	.dataa(!\D_iw[16]~q ),
	.datab(!\D_iw[12]~q ),
	.datac(!\D_iw[11]~q ),
	.datad(!\Equal4~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_jmp_indirect~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_jmp_indirect~0 .extended_lut = "off";
defparam \D_ctrl_jmp_indirect~0 .lut_mask = 64'hEFFFEFFFEFFFEFFF;
defparam \D_ctrl_jmp_indirect~0 .shared_arith = "off";

dffeas E_ctrl_jmp_indirect(
	.clk(clk_clk),
	.d(\D_ctrl_jmp_indirect~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_ctrl_jmp_indirect~q ),
	.prn(vcc));
defparam E_ctrl_jmp_indirect.is_wysiwyg = "true";
defparam E_ctrl_jmp_indirect.power_up = "low";

dffeas E_ctrl_jmp_direct(
	.clk(clk_clk),
	.d(\D_ctrl_a_not_src~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_ctrl_jmp_direct~q ),
	.prn(vcc));
defparam E_ctrl_jmp_direct.is_wysiwyg = "true";
defparam E_ctrl_jmp_direct.power_up = "low";

cyclonev_lcell_comb \M_pipe_flush_waddr[7]~0 (
	.dataa(!\E_ctrl_break~q ),
	.datab(!\E_ctrl_exception~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_pipe_flush_waddr[7]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_pipe_flush_waddr[7]~0 .extended_lut = "off";
defparam \M_pipe_flush_waddr[7]~0 .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \M_pipe_flush_waddr[7]~0 .shared_arith = "off";

cyclonev_lcell_comb \Add3~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\F_pc[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add3~57_sumout ),
	.cout(\Add3~58 ),
	.shareout());
defparam \Add3~57 .extended_lut = "off";
defparam \Add3~57 .lut_mask = 64'h00000000000000FF;
defparam \Add3~57 .shared_arith = "off";

cyclonev_lcell_comb \Add0~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\processor_cpu_ic_data|the_altsyncram|auto_generated|q_b[8] ),
	.datae(gnd),
	.dataf(!\Add3~57_sumout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~37_sumout ),
	.cout(\Add0~38 ),
	.shareout());
defparam \Add0~37 .extended_lut = "off";
defparam \Add0~37 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~37 .shared_arith = "off";

dffeas \D_br_taken_waddr_partial[0] (
	.clk(clk_clk),
	.d(\Add0~37_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\D_br_taken_waddr_partial[0]~q ),
	.prn(vcc));
defparam \D_br_taken_waddr_partial[0] .is_wysiwyg = "true";
defparam \D_br_taken_waddr_partial[0] .power_up = "low";

dffeas \D_pc_plus_one[0] (
	.clk(clk_clk),
	.d(\Add3~57_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\D_pc_plus_one[0]~q ),
	.prn(vcc));
defparam \D_pc_plus_one[0] .is_wysiwyg = "true";
defparam \D_pc_plus_one[0] .power_up = "low";

cyclonev_lcell_comb D_br_pred_not_taken(
	.dataa(!\D_iw[0]~q ),
	.datab(!\D_iw[1]~q ),
	.datac(!\D_iw[21]~q ),
	.datad(!\E_ctrl_br_cond_nxt~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_br_pred_not_taken~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam D_br_pred_not_taken.extended_lut = "off";
defparam D_br_pred_not_taken.lut_mask = 64'hDFFFDFFFDFFFDFFF;
defparam D_br_pred_not_taken.shared_arith = "off";

dffeas \E_extra_pc[0] (
	.clk(clk_clk),
	.d(\D_br_taken_waddr_partial[0]~q ),
	.asdata(\D_pc_plus_one[0]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\D_br_pred_not_taken~combout ),
	.ena(\W_stall~combout ),
	.q(\E_extra_pc[0]~q ),
	.prn(vcc));
defparam \E_extra_pc[0] .is_wysiwyg = "true";
defparam \E_extra_pc[0] .power_up = "low";

cyclonev_lcell_comb \M_pipe_flush_waddr[7]~1 (
	.dataa(!\E_ctrl_jmp_indirect~q ),
	.datab(!\E_ctrl_jmp_direct~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_pipe_flush_waddr[7]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_pipe_flush_waddr[7]~1 .extended_lut = "off";
defparam \M_pipe_flush_waddr[7]~1 .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \M_pipe_flush_waddr[7]~1 .shared_arith = "off";

cyclonev_lcell_comb \M_pipe_flush_waddr_nxt[0]~0 (
	.dataa(!\E_src1[2]~24_combout ),
	.datab(!\E_src1[2]~25_combout ),
	.datac(!\E_extra_pc[0]~q ),
	.datad(!\M_pipe_flush_waddr[7]~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_pipe_flush_waddr_nxt[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_pipe_flush_waddr_nxt[0]~0 .extended_lut = "off";
defparam \M_pipe_flush_waddr_nxt[0]~0 .lut_mask = 64'hFAFCFAFCFAFCFAFC;
defparam \M_pipe_flush_waddr_nxt[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \M_pipe_flush_waddr_nxt[0]~1 (
	.dataa(!\E_hbreak_req~combout ),
	.datab(!\E_iw[6]~q ),
	.datac(!\E_ctrl_jmp_indirect~q ),
	.datad(!\E_ctrl_jmp_direct~q ),
	.datae(!\M_pipe_flush_waddr[7]~0_combout ),
	.dataf(!\M_pipe_flush_waddr_nxt[0]~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_pipe_flush_waddr_nxt[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_pipe_flush_waddr_nxt[0]~1 .extended_lut = "off";
defparam \M_pipe_flush_waddr_nxt[0]~1 .lut_mask = 64'hFFFFFFFF7FF7FFFF;
defparam \M_pipe_flush_waddr_nxt[0]~1 .shared_arith = "off";

dffeas \D_pc[0] (
	.clk(clk_clk),
	.d(\F_pc[0]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\D_pc[0]~q ),
	.prn(vcc));
defparam \D_pc[0] .is_wysiwyg = "true";
defparam \D_pc[0] .power_up = "low";

dffeas \E_pc[0] (
	.clk(clk_clk),
	.d(\D_pc[0]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_pc[0]~q ),
	.prn(vcc));
defparam \E_pc[0] .is_wysiwyg = "true";
defparam \E_pc[0] .power_up = "low";

cyclonev_lcell_comb \M_pipe_flush_waddr[7]~2 (
	.dataa(!\E_hbreak_req~combout ),
	.datab(!\E_ctrl_crst~q ),
	.datac(!\M_pipe_flush_waddr[7]~1_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_pipe_flush_waddr[7]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_pipe_flush_waddr[7]~2 .extended_lut = "off";
defparam \M_pipe_flush_waddr[7]~2 .lut_mask = 64'hBFBFBFBFBFBFBFBF;
defparam \M_pipe_flush_waddr[7]~2 .shared_arith = "off";

dffeas \M_pipe_flush_waddr[0] (
	.clk(clk_clk),
	.d(\M_pipe_flush_waddr_nxt[0]~1_combout ),
	.asdata(\E_pc[0]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\M_pipe_flush_waddr[7]~2_combout ),
	.sload(\E_hbreak_req~combout ),
	.ena(\W_stall~combout ),
	.q(\M_pipe_flush_waddr[0]~q ),
	.prn(vcc));
defparam \M_pipe_flush_waddr[0] .is_wysiwyg = "true";
defparam \M_pipe_flush_waddr[0] .power_up = "low";

cyclonev_lcell_comb \F_ic_data_rd_addr_nxt[0]~0 (
	.dataa(!\M_pipe_flush~q ),
	.datab(!\D_iw[21]~q ),
	.datac(!\D_issue~q ),
	.datad(!\D_ctrl_br~0_combout ),
	.datae(!\D_refetch~0_combout ),
	.dataf(!\Equal4~12_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ic_data_rd_addr_nxt[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ic_data_rd_addr_nxt[0]~0 .extended_lut = "off";
defparam \F_ic_data_rd_addr_nxt[0]~0 .lut_mask = 64'h7FFFFFFFFFFFFFFF;
defparam \F_ic_data_rd_addr_nxt[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \F_ic_data_rd_addr_nxt[0]~1 (
	.dataa(!\M_pipe_flush_waddr[0]~q ),
	.datab(!\D_pc[0]~q ),
	.datac(!\Add3~57_sumout ),
	.datad(!\D_br_taken_waddr_partial[0]~q ),
	.datae(!\F_ic_data_rd_addr_nxt[0]~0_combout ),
	.dataf(!\F_kill~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ic_data_rd_addr_nxt[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ic_data_rd_addr_nxt[0]~1 .extended_lut = "off";
defparam \F_ic_data_rd_addr_nxt[0]~1 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \F_ic_data_rd_addr_nxt[0]~1 .shared_arith = "off";

dffeas \F_pc[0] (
	.clk(clk_clk),
	.d(\F_ic_data_rd_addr_nxt[0]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\F_pc[0]~q ),
	.prn(vcc));
defparam \F_pc[0] .is_wysiwyg = "true";
defparam \F_pc[0] .power_up = "low";

cyclonev_lcell_comb \Add3~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\F_pc[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~58 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add3~53_sumout ),
	.cout(\Add3~54 ),
	.shareout());
defparam \Add3~53 .extended_lut = "off";
defparam \Add3~53 .lut_mask = 64'h00000000000000FF;
defparam \Add3~53 .shared_arith = "off";

cyclonev_lcell_comb \Add0~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\processor_cpu_ic_data|the_altsyncram|auto_generated|q_b[9] ),
	.datae(gnd),
	.dataf(!\Add3~53_sumout ),
	.datag(gnd),
	.cin(\Add0~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~33_sumout ),
	.cout(\Add0~34 ),
	.shareout());
defparam \Add0~33 .extended_lut = "off";
defparam \Add0~33 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~33 .shared_arith = "off";

dffeas \D_br_taken_waddr_partial[1] (
	.clk(clk_clk),
	.d(\Add0~33_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\D_br_taken_waddr_partial[1]~q ),
	.prn(vcc));
defparam \D_br_taken_waddr_partial[1] .is_wysiwyg = "true";
defparam \D_br_taken_waddr_partial[1] .power_up = "low";

dffeas \D_pc_plus_one[1] (
	.clk(clk_clk),
	.d(\Add3~53_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\D_pc_plus_one[1]~q ),
	.prn(vcc));
defparam \D_pc_plus_one[1] .is_wysiwyg = "true";
defparam \D_pc_plus_one[1] .power_up = "low";

dffeas \E_extra_pc[1] (
	.clk(clk_clk),
	.d(\D_br_taken_waddr_partial[1]~q ),
	.asdata(\D_pc_plus_one[1]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\D_br_pred_not_taken~combout ),
	.ena(\W_stall~combout ),
	.q(\E_extra_pc[1]~q ),
	.prn(vcc));
defparam \E_extra_pc[1] .is_wysiwyg = "true";
defparam \E_extra_pc[1] .power_up = "low";

cyclonev_lcell_comb \M_pipe_flush_waddr_nxt[1]~2 (
	.dataa(!\E_extra_pc[1]~q ),
	.datab(!\M_wr_data_unfiltered[3]~8_combout ),
	.datac(!\E_src1_hazard_M~q ),
	.datad(!\E_src1_prelim[3]~q ),
	.datae(!\M_pipe_flush_waddr[7]~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_pipe_flush_waddr_nxt[1]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_pipe_flush_waddr_nxt[1]~2 .extended_lut = "off";
defparam \M_pipe_flush_waddr_nxt[1]~2 .lut_mask = 64'h7FFFF7FF7FFFF7FF;
defparam \M_pipe_flush_waddr_nxt[1]~2 .shared_arith = "off";

cyclonev_lcell_comb \M_pipe_flush_waddr_nxt[1]~3 (
	.dataa(!\E_hbreak_req~combout ),
	.datab(!\E_iw[7]~q ),
	.datac(!\E_ctrl_jmp_indirect~q ),
	.datad(!\E_ctrl_jmp_direct~q ),
	.datae(!\M_pipe_flush_waddr[7]~0_combout ),
	.dataf(!\M_pipe_flush_waddr_nxt[1]~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_pipe_flush_waddr_nxt[1]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_pipe_flush_waddr_nxt[1]~3 .extended_lut = "off";
defparam \M_pipe_flush_waddr_nxt[1]~3 .lut_mask = 64'h7FF7FFFFFFFFFFFF;
defparam \M_pipe_flush_waddr_nxt[1]~3 .shared_arith = "off";

dffeas \D_pc[1] (
	.clk(clk_clk),
	.d(\F_pc[1]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\D_pc[1]~q ),
	.prn(vcc));
defparam \D_pc[1] .is_wysiwyg = "true";
defparam \D_pc[1] .power_up = "low";

dffeas \E_pc[1] (
	.clk(clk_clk),
	.d(\D_pc[1]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_pc[1]~q ),
	.prn(vcc));
defparam \E_pc[1] .is_wysiwyg = "true";
defparam \E_pc[1] .power_up = "low";

dffeas \M_pipe_flush_waddr[1] (
	.clk(clk_clk),
	.d(\M_pipe_flush_waddr_nxt[1]~3_combout ),
	.asdata(\E_pc[1]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\M_pipe_flush_waddr[7]~2_combout ),
	.sload(\E_hbreak_req~combout ),
	.ena(\W_stall~combout ),
	.q(\M_pipe_flush_waddr[1]~q ),
	.prn(vcc));
defparam \M_pipe_flush_waddr[1] .is_wysiwyg = "true";
defparam \M_pipe_flush_waddr[1] .power_up = "low";

cyclonev_lcell_comb \F_ic_data_rd_addr_nxt[1]~2 (
	.dataa(!\M_pipe_flush_waddr[1]~q ),
	.datab(!\D_pc[1]~q ),
	.datac(!\Add3~53_sumout ),
	.datad(!\D_br_taken_waddr_partial[1]~q ),
	.datae(!\F_ic_data_rd_addr_nxt[0]~0_combout ),
	.dataf(!\F_kill~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ic_data_rd_addr_nxt[1]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ic_data_rd_addr_nxt[1]~2 .extended_lut = "off";
defparam \F_ic_data_rd_addr_nxt[1]~2 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \F_ic_data_rd_addr_nxt[1]~2 .shared_arith = "off";

dffeas \F_pc[1] (
	.clk(clk_clk),
	.d(\F_ic_data_rd_addr_nxt[1]~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\F_pc[1]~q ),
	.prn(vcc));
defparam \F_pc[1] .is_wysiwyg = "true";
defparam \F_pc[1] .power_up = "low";

cyclonev_lcell_comb \Add3~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\F_pc[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~54 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add3~5_sumout ),
	.cout(\Add3~6 ),
	.shareout());
defparam \Add3~5 .extended_lut = "off";
defparam \Add3~5 .lut_mask = 64'h00000000000000FF;
defparam \Add3~5 .shared_arith = "off";

cyclonev_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\processor_cpu_ic_data|the_altsyncram|auto_generated|q_b[10] ),
	.datae(gnd),
	.dataf(!\Add3~5_sumout ),
	.datag(gnd),
	.cin(\Add0~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout());
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~5 .shared_arith = "off";

dffeas \D_br_taken_waddr_partial[2] (
	.clk(clk_clk),
	.d(\Add0~5_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\D_br_taken_waddr_partial[2]~q ),
	.prn(vcc));
defparam \D_br_taken_waddr_partial[2] .is_wysiwyg = "true";
defparam \D_br_taken_waddr_partial[2] .power_up = "low";

dffeas \D_pc_plus_one[2] (
	.clk(clk_clk),
	.d(\Add3~5_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\D_pc_plus_one[2]~q ),
	.prn(vcc));
defparam \D_pc_plus_one[2] .is_wysiwyg = "true";
defparam \D_pc_plus_one[2] .power_up = "low";

dffeas \E_extra_pc[2] (
	.clk(clk_clk),
	.d(\D_br_taken_waddr_partial[2]~q ),
	.asdata(\D_pc_plus_one[2]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\D_br_pred_not_taken~combout ),
	.ena(\W_stall~combout ),
	.q(\E_extra_pc[2]~q ),
	.prn(vcc));
defparam \E_extra_pc[2] .is_wysiwyg = "true";
defparam \E_extra_pc[2] .power_up = "low";

cyclonev_lcell_comb \M_pipe_flush_waddr_nxt[2]~4 (
	.dataa(!\E_src1[4]~1_combout ),
	.datab(!\E_src1[4]~2_combout ),
	.datac(!\E_extra_pc[2]~q ),
	.datad(!\M_pipe_flush_waddr[7]~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_pipe_flush_waddr_nxt[2]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_pipe_flush_waddr_nxt[2]~4 .extended_lut = "off";
defparam \M_pipe_flush_waddr_nxt[2]~4 .lut_mask = 64'hFAFCFAFCFAFCFAFC;
defparam \M_pipe_flush_waddr_nxt[2]~4 .shared_arith = "off";

cyclonev_lcell_comb \M_pipe_flush_waddr_nxt[2]~5 (
	.dataa(!\E_hbreak_req~combout ),
	.datab(!\E_iw[8]~q ),
	.datac(!\E_ctrl_jmp_indirect~q ),
	.datad(!\E_ctrl_jmp_direct~q ),
	.datae(!\M_pipe_flush_waddr[7]~0_combout ),
	.dataf(!\M_pipe_flush_waddr_nxt[2]~4_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_pipe_flush_waddr_nxt[2]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_pipe_flush_waddr_nxt[2]~5 .extended_lut = "off";
defparam \M_pipe_flush_waddr_nxt[2]~5 .lut_mask = 64'hFFFFFFFF7FF7FFFF;
defparam \M_pipe_flush_waddr_nxt[2]~5 .shared_arith = "off";

dffeas \D_pc[2] (
	.clk(clk_clk),
	.d(\F_pc[2]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\D_pc[2]~q ),
	.prn(vcc));
defparam \D_pc[2] .is_wysiwyg = "true";
defparam \D_pc[2] .power_up = "low";

dffeas \E_pc[2] (
	.clk(clk_clk),
	.d(\D_pc[2]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_pc[2]~q ),
	.prn(vcc));
defparam \E_pc[2] .is_wysiwyg = "true";
defparam \E_pc[2] .power_up = "low";

dffeas \M_pipe_flush_waddr[2] (
	.clk(clk_clk),
	.d(\M_pipe_flush_waddr_nxt[2]~5_combout ),
	.asdata(\E_pc[2]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\M_pipe_flush_waddr[7]~2_combout ),
	.sload(\E_hbreak_req~combout ),
	.ena(\W_stall~combout ),
	.q(\M_pipe_flush_waddr[2]~q ),
	.prn(vcc));
defparam \M_pipe_flush_waddr[2] .is_wysiwyg = "true";
defparam \M_pipe_flush_waddr[2] .power_up = "low";

cyclonev_lcell_comb \F_ic_data_rd_addr_nxt[2]~3 (
	.dataa(!\M_pipe_flush_waddr[2]~q ),
	.datab(!\D_pc[2]~q ),
	.datac(!\Add3~5_sumout ),
	.datad(!\D_br_taken_waddr_partial[2]~q ),
	.datae(!\F_ic_data_rd_addr_nxt[0]~0_combout ),
	.dataf(!\F_kill~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ic_data_rd_addr_nxt[2]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ic_data_rd_addr_nxt[2]~3 .extended_lut = "off";
defparam \F_ic_data_rd_addr_nxt[2]~3 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \F_ic_data_rd_addr_nxt[2]~3 .shared_arith = "off";

dffeas \F_pc[2] (
	.clk(clk_clk),
	.d(\F_ic_data_rd_addr_nxt[2]~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\F_pc[2]~q ),
	.prn(vcc));
defparam \F_pc[2] .is_wysiwyg = "true";
defparam \F_pc[2] .power_up = "low";

cyclonev_lcell_comb \F_ic_valid~4 (
	.dataa(!\processor_cpu_ic_tag|the_altsyncram|auto_generated|q_b[7] ),
	.datab(!\processor_cpu_ic_tag|the_altsyncram|auto_generated|q_b[9] ),
	.datac(!\processor_cpu_ic_tag|the_altsyncram|auto_generated|q_b[8] ),
	.datad(!\F_pc[0]~q ),
	.datae(!\F_pc[1]~q ),
	.dataf(!\F_pc[2]~q ),
	.datag(!\processor_cpu_ic_tag|the_altsyncram|auto_generated|q_b[6] ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ic_valid~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ic_valid~4 .extended_lut = "on";
defparam \F_ic_valid~4 .lut_mask = 64'hFAFCFAFCFAFCFAFC;
defparam \F_ic_valid~4 .shared_arith = "off";

cyclonev_lcell_comb \F_ic_valid~0 (
	.dataa(!\processor_cpu_ic_tag|the_altsyncram|auto_generated|q_b[11] ),
	.datab(!\processor_cpu_ic_tag|the_altsyncram|auto_generated|q_b[13] ),
	.datac(!\processor_cpu_ic_tag|the_altsyncram|auto_generated|q_b[12] ),
	.datad(!\F_pc[2]~q ),
	.datae(!\F_pc[1]~q ),
	.dataf(!\F_ic_valid~4_combout ),
	.datag(!\processor_cpu_ic_tag|the_altsyncram|auto_generated|q_b[10] ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ic_valid~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ic_valid~0 .extended_lut = "on";
defparam \F_ic_valid~0 .lut_mask = 64'hFAFCFAFCFAFCFAFC;
defparam \F_ic_valid~0 .shared_arith = "off";

dffeas \D_pc[13] (
	.clk(clk_clk),
	.d(\F_pc[13]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\D_pc[13]~q ),
	.prn(vcc));
defparam \D_pc[13] .is_wysiwyg = "true";
defparam \D_pc[13] .power_up = "low";

dffeas \E_pc[13] (
	.clk(clk_clk),
	.d(\D_pc[13]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_pc[13]~q ),
	.prn(vcc));
defparam \E_pc[13] .is_wysiwyg = "true";
defparam \E_pc[13] .power_up = "low";

cyclonev_lcell_comb \Add3~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\F_pc[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add3~1_sumout ),
	.cout(\Add3~2 ),
	.shareout());
defparam \Add3~1 .extended_lut = "off";
defparam \Add3~1 .lut_mask = 64'h00000000000000FF;
defparam \Add3~1 .shared_arith = "off";

cyclonev_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\processor_cpu_ic_data|the_altsyncram|auto_generated|q_b[11] ),
	.datae(gnd),
	.dataf(!\Add3~1_sumout ),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(\Add0~2 ),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~1 .shared_arith = "off";

dffeas \D_br_taken_waddr_partial[3] (
	.clk(clk_clk),
	.d(\Add0~1_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\D_br_taken_waddr_partial[3]~q ),
	.prn(vcc));
defparam \D_br_taken_waddr_partial[3] .is_wysiwyg = "true";
defparam \D_br_taken_waddr_partial[3] .power_up = "low";

dffeas \D_pc_plus_one[3] (
	.clk(clk_clk),
	.d(\Add3~1_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\D_pc_plus_one[3]~q ),
	.prn(vcc));
defparam \D_pc_plus_one[3] .is_wysiwyg = "true";
defparam \D_pc_plus_one[3] .power_up = "low";

dffeas \E_extra_pc[3] (
	.clk(clk_clk),
	.d(\D_br_taken_waddr_partial[3]~q ),
	.asdata(\D_pc_plus_one[3]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\D_br_pred_not_taken~combout ),
	.ena(\W_stall~combout ),
	.q(\E_extra_pc[3]~q ),
	.prn(vcc));
defparam \E_extra_pc[3] .is_wysiwyg = "true";
defparam \E_extra_pc[3] .power_up = "low";

cyclonev_lcell_comb \M_pipe_flush_waddr_nxt[3]~6 (
	.dataa(!\E_src1_hazard_M~q ),
	.datab(!\E_extra_pc[3]~q ),
	.datac(!\M_wr_data_unfiltered[5]~0_combout ),
	.datad(!\E_src1_prelim[5]~q ),
	.datae(!\M_pipe_flush_waddr[7]~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_pipe_flush_waddr_nxt[3]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_pipe_flush_waddr_nxt[3]~6 .extended_lut = "off";
defparam \M_pipe_flush_waddr_nxt[3]~6 .lut_mask = 64'h7FFFBFFF7FFFBFFF;
defparam \M_pipe_flush_waddr_nxt[3]~6 .shared_arith = "off";

dffeas \E_iw[9] (
	.clk(clk_clk),
	.d(\D_iw[9]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_iw[9]~q ),
	.prn(vcc));
defparam \E_iw[9] .is_wysiwyg = "true";
defparam \E_iw[9] .power_up = "low";

cyclonev_lcell_comb \M_pipe_flush_waddr_nxt[3]~7 (
	.dataa(!\E_hbreak_req~combout ),
	.datab(!\E_ctrl_jmp_indirect~q ),
	.datac(!\E_ctrl_jmp_direct~q ),
	.datad(!\M_pipe_flush_waddr[7]~0_combout ),
	.datae(!\M_pipe_flush_waddr_nxt[3]~6_combout ),
	.dataf(!\E_iw[9]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_pipe_flush_waddr_nxt[3]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_pipe_flush_waddr_nxt[3]~7 .extended_lut = "off";
defparam \M_pipe_flush_waddr_nxt[3]~7 .lut_mask = 64'hFFBEFFFFFFFFFFFF;
defparam \M_pipe_flush_waddr_nxt[3]~7 .shared_arith = "off";

dffeas \D_pc[3] (
	.clk(clk_clk),
	.d(\F_pc[3]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\D_pc[3]~q ),
	.prn(vcc));
defparam \D_pc[3] .is_wysiwyg = "true";
defparam \D_pc[3] .power_up = "low";

dffeas \E_pc[3] (
	.clk(clk_clk),
	.d(\D_pc[3]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_pc[3]~q ),
	.prn(vcc));
defparam \E_pc[3] .is_wysiwyg = "true";
defparam \E_pc[3] .power_up = "low";

dffeas \M_pipe_flush_waddr[3] (
	.clk(clk_clk),
	.d(\M_pipe_flush_waddr_nxt[3]~7_combout ),
	.asdata(\E_pc[3]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\M_pipe_flush_waddr[7]~2_combout ),
	.sload(\E_hbreak_req~combout ),
	.ena(\W_stall~combout ),
	.q(\M_pipe_flush_waddr[3]~q ),
	.prn(vcc));
defparam \M_pipe_flush_waddr[3] .is_wysiwyg = "true";
defparam \M_pipe_flush_waddr[3] .power_up = "low";

cyclonev_lcell_comb \F_ic_tag_rd_addr_nxt[0]~0 (
	.dataa(!\M_pipe_flush_waddr[3]~q ),
	.datab(!\D_pc[3]~q ),
	.datac(!\Add3~1_sumout ),
	.datad(!\D_br_taken_waddr_partial[3]~q ),
	.datae(!\F_ic_data_rd_addr_nxt[0]~0_combout ),
	.dataf(!\F_kill~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ic_tag_rd_addr_nxt[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ic_tag_rd_addr_nxt[0]~0 .extended_lut = "off";
defparam \F_ic_tag_rd_addr_nxt[0]~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \F_ic_tag_rd_addr_nxt[0]~0 .shared_arith = "off";

dffeas \F_pc[3] (
	.clk(clk_clk),
	.d(\F_ic_tag_rd_addr_nxt[0]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\F_pc[3]~q ),
	.prn(vcc));
defparam \F_pc[3] .is_wysiwyg = "true";
defparam \F_pc[3] .power_up = "low";

cyclonev_lcell_comb \Add3~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\F_pc[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add3~9_sumout ),
	.cout(\Add3~10 ),
	.shareout());
defparam \Add3~9 .extended_lut = "off";
defparam \Add3~9 .lut_mask = 64'h00000000000000FF;
defparam \Add3~9 .shared_arith = "off";

cyclonev_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\processor_cpu_ic_data|the_altsyncram|auto_generated|q_b[12] ),
	.datae(gnd),
	.dataf(!\Add3~9_sumout ),
	.datag(gnd),
	.cin(\Add0~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout());
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~9 .shared_arith = "off";

dffeas \D_br_taken_waddr_partial[4] (
	.clk(clk_clk),
	.d(\Add0~9_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\D_br_taken_waddr_partial[4]~q ),
	.prn(vcc));
defparam \D_br_taken_waddr_partial[4] .is_wysiwyg = "true";
defparam \D_br_taken_waddr_partial[4] .power_up = "low";

dffeas \D_pc_plus_one[4] (
	.clk(clk_clk),
	.d(\Add3~9_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\D_pc_plus_one[4]~q ),
	.prn(vcc));
defparam \D_pc_plus_one[4] .is_wysiwyg = "true";
defparam \D_pc_plus_one[4] .power_up = "low";

dffeas \E_extra_pc[4] (
	.clk(clk_clk),
	.d(\D_br_taken_waddr_partial[4]~q ),
	.asdata(\D_pc_plus_one[4]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\D_br_pred_not_taken~combout ),
	.ena(\W_stall~combout ),
	.q(\E_extra_pc[4]~q ),
	.prn(vcc));
defparam \E_extra_pc[4] .is_wysiwyg = "true";
defparam \E_extra_pc[4] .power_up = "low";

cyclonev_lcell_comb \M_pipe_flush_waddr_nxt[4]~8 (
	.dataa(!\E_extra_pc[4]~q ),
	.datab(!\E_src1[6]~4_combout ),
	.datac(!\E_src1[6]~5_combout ),
	.datad(!\M_pipe_flush_waddr[7]~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_pipe_flush_waddr_nxt[4]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_pipe_flush_waddr_nxt[4]~8 .extended_lut = "off";
defparam \M_pipe_flush_waddr_nxt[4]~8 .lut_mask = 64'hFAFCFAFCFAFCFAFC;
defparam \M_pipe_flush_waddr_nxt[4]~8 .shared_arith = "off";

dffeas \E_iw[10] (
	.clk(clk_clk),
	.d(\D_iw[10]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_iw[10]~q ),
	.prn(vcc));
defparam \E_iw[10] .is_wysiwyg = "true";
defparam \E_iw[10] .power_up = "low";

cyclonev_lcell_comb \M_pipe_flush_waddr_nxt[4]~9 (
	.dataa(!\E_hbreak_req~combout ),
	.datab(!\E_ctrl_jmp_indirect~q ),
	.datac(!\E_ctrl_jmp_direct~q ),
	.datad(!\M_pipe_flush_waddr[7]~0_combout ),
	.datae(!\M_pipe_flush_waddr_nxt[4]~8_combout ),
	.dataf(!\E_iw[10]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_pipe_flush_waddr_nxt[4]~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_pipe_flush_waddr_nxt[4]~9 .extended_lut = "off";
defparam \M_pipe_flush_waddr_nxt[4]~9 .lut_mask = 64'hFFFF7DFFFFFFFFFF;
defparam \M_pipe_flush_waddr_nxt[4]~9 .shared_arith = "off";

dffeas \D_pc[4] (
	.clk(clk_clk),
	.d(\F_pc[4]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\D_pc[4]~q ),
	.prn(vcc));
defparam \D_pc[4] .is_wysiwyg = "true";
defparam \D_pc[4] .power_up = "low";

dffeas \E_pc[4] (
	.clk(clk_clk),
	.d(\D_pc[4]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_pc[4]~q ),
	.prn(vcc));
defparam \E_pc[4] .is_wysiwyg = "true";
defparam \E_pc[4] .power_up = "low";

dffeas \M_pipe_flush_waddr[4] (
	.clk(clk_clk),
	.d(\M_pipe_flush_waddr_nxt[4]~9_combout ),
	.asdata(\E_pc[4]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\M_pipe_flush_waddr[7]~2_combout ),
	.sload(\E_hbreak_req~combout ),
	.ena(\W_stall~combout ),
	.q(\M_pipe_flush_waddr[4]~q ),
	.prn(vcc));
defparam \M_pipe_flush_waddr[4] .is_wysiwyg = "true";
defparam \M_pipe_flush_waddr[4] .power_up = "low";

cyclonev_lcell_comb \F_ic_tag_rd_addr_nxt[1]~1 (
	.dataa(!\M_pipe_flush_waddr[4]~q ),
	.datab(!\D_pc[4]~q ),
	.datac(!\Add3~9_sumout ),
	.datad(!\D_br_taken_waddr_partial[4]~q ),
	.datae(!\F_ic_data_rd_addr_nxt[0]~0_combout ),
	.dataf(!\F_kill~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ic_tag_rd_addr_nxt[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ic_tag_rd_addr_nxt[1]~1 .extended_lut = "off";
defparam \F_ic_tag_rd_addr_nxt[1]~1 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \F_ic_tag_rd_addr_nxt[1]~1 .shared_arith = "off";

dffeas \F_pc[4] (
	.clk(clk_clk),
	.d(\F_ic_tag_rd_addr_nxt[1]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\F_pc[4]~q ),
	.prn(vcc));
defparam \F_pc[4] .is_wysiwyg = "true";
defparam \F_pc[4] .power_up = "low";

cyclonev_lcell_comb \Add3~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\F_pc[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add3~49_sumout ),
	.cout(\Add3~50 ),
	.shareout());
defparam \Add3~49 .extended_lut = "off";
defparam \Add3~49 .lut_mask = 64'h00000000000000FF;
defparam \Add3~49 .shared_arith = "off";

cyclonev_lcell_comb \Add0~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\processor_cpu_ic_data|the_altsyncram|auto_generated|q_b[13] ),
	.datae(gnd),
	.dataf(!\Add3~49_sumout ),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~29_sumout ),
	.cout(\Add0~30 ),
	.shareout());
defparam \Add0~29 .extended_lut = "off";
defparam \Add0~29 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~29 .shared_arith = "off";

dffeas \D_br_taken_waddr_partial[5] (
	.clk(clk_clk),
	.d(\Add0~29_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\D_br_taken_waddr_partial[5]~q ),
	.prn(vcc));
defparam \D_br_taken_waddr_partial[5] .is_wysiwyg = "true";
defparam \D_br_taken_waddr_partial[5] .power_up = "low";

dffeas \D_pc_plus_one[5] (
	.clk(clk_clk),
	.d(\Add3~49_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\D_pc_plus_one[5]~q ),
	.prn(vcc));
defparam \D_pc_plus_one[5] .is_wysiwyg = "true";
defparam \D_pc_plus_one[5] .power_up = "low";

dffeas \E_extra_pc[5] (
	.clk(clk_clk),
	.d(\D_br_taken_waddr_partial[5]~q ),
	.asdata(\D_pc_plus_one[5]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\D_br_pred_not_taken~combout ),
	.ena(\W_stall~combout ),
	.q(\E_extra_pc[5]~q ),
	.prn(vcc));
defparam \E_extra_pc[5] .is_wysiwyg = "true";
defparam \E_extra_pc[5] .power_up = "low";

cyclonev_lcell_comb \M_pipe_flush_waddr_nxt[5]~10 (
	.dataa(!\E_src1_hazard_M~q ),
	.datab(!\M_wr_data_unfiltered[7]~7_combout ),
	.datac(!\E_src1_prelim[7]~q ),
	.datad(!\E_extra_pc[5]~q ),
	.datae(!\M_pipe_flush_waddr[7]~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_pipe_flush_waddr_nxt[5]~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_pipe_flush_waddr_nxt[5]~10 .extended_lut = "off";
defparam \M_pipe_flush_waddr_nxt[5]~10 .lut_mask = 64'h7FFFBFFF7FFFBFFF;
defparam \M_pipe_flush_waddr_nxt[5]~10 .shared_arith = "off";

cyclonev_lcell_comb \M_pipe_flush_waddr_nxt[5]~11 (
	.dataa(!\E_iw[11]~q ),
	.datab(!\E_hbreak_req~combout ),
	.datac(!\E_ctrl_jmp_indirect~q ),
	.datad(!\E_ctrl_jmp_direct~q ),
	.datae(!\M_pipe_flush_waddr[7]~0_combout ),
	.dataf(!\M_pipe_flush_waddr_nxt[5]~10_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_pipe_flush_waddr_nxt[5]~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_pipe_flush_waddr_nxt[5]~11 .extended_lut = "off";
defparam \M_pipe_flush_waddr_nxt[5]~11 .lut_mask = 64'h7FF7FFFFFFFFFFFF;
defparam \M_pipe_flush_waddr_nxt[5]~11 .shared_arith = "off";

dffeas \D_pc[5] (
	.clk(clk_clk),
	.d(\F_pc[5]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\D_pc[5]~q ),
	.prn(vcc));
defparam \D_pc[5] .is_wysiwyg = "true";
defparam \D_pc[5] .power_up = "low";

dffeas \E_pc[5] (
	.clk(clk_clk),
	.d(\D_pc[5]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_pc[5]~q ),
	.prn(vcc));
defparam \E_pc[5] .is_wysiwyg = "true";
defparam \E_pc[5] .power_up = "low";

dffeas \M_pipe_flush_waddr[5] (
	.clk(clk_clk),
	.d(\M_pipe_flush_waddr_nxt[5]~11_combout ),
	.asdata(\E_pc[5]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\M_pipe_flush_waddr[7]~2_combout ),
	.sload(\E_hbreak_req~combout ),
	.ena(\W_stall~combout ),
	.q(\M_pipe_flush_waddr[5]~q ),
	.prn(vcc));
defparam \M_pipe_flush_waddr[5] .is_wysiwyg = "true";
defparam \M_pipe_flush_waddr[5] .power_up = "low";

cyclonev_lcell_comb \F_ic_tag_rd_addr_nxt[2]~2 (
	.dataa(!\M_pipe_flush_waddr[5]~q ),
	.datab(!\D_pc[5]~q ),
	.datac(!\Add3~49_sumout ),
	.datad(!\D_br_taken_waddr_partial[5]~q ),
	.datae(!\F_ic_data_rd_addr_nxt[0]~0_combout ),
	.dataf(!\F_kill~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ic_tag_rd_addr_nxt[2]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ic_tag_rd_addr_nxt[2]~2 .extended_lut = "off";
defparam \F_ic_tag_rd_addr_nxt[2]~2 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \F_ic_tag_rd_addr_nxt[2]~2 .shared_arith = "off";

dffeas \F_pc[5] (
	.clk(clk_clk),
	.d(\F_ic_tag_rd_addr_nxt[2]~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\F_pc[5]~q ),
	.prn(vcc));
defparam \F_pc[5] .is_wysiwyg = "true";
defparam \F_pc[5] .power_up = "low";

cyclonev_lcell_comb \Add3~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\F_pc[6]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~50 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add3~45_sumout ),
	.cout(\Add3~46 ),
	.shareout());
defparam \Add3~45 .extended_lut = "off";
defparam \Add3~45 .lut_mask = 64'h00000000000000FF;
defparam \Add3~45 .shared_arith = "off";

cyclonev_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\processor_cpu_ic_data|the_altsyncram|auto_generated|q_b[14] ),
	.datae(gnd),
	.dataf(!\Add3~45_sumout ),
	.datag(gnd),
	.cin(\Add0~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout());
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~25 .shared_arith = "off";

dffeas \D_br_taken_waddr_partial[6] (
	.clk(clk_clk),
	.d(\Add0~25_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\D_br_taken_waddr_partial[6]~q ),
	.prn(vcc));
defparam \D_br_taken_waddr_partial[6] .is_wysiwyg = "true";
defparam \D_br_taken_waddr_partial[6] .power_up = "low";

dffeas \D_pc_plus_one[6] (
	.clk(clk_clk),
	.d(\Add3~45_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\D_pc_plus_one[6]~q ),
	.prn(vcc));
defparam \D_pc_plus_one[6] .is_wysiwyg = "true";
defparam \D_pc_plus_one[6] .power_up = "low";

dffeas \E_extra_pc[6] (
	.clk(clk_clk),
	.d(\D_br_taken_waddr_partial[6]~q ),
	.asdata(\D_pc_plus_one[6]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\D_br_pred_not_taken~combout ),
	.ena(\W_stall~combout ),
	.q(\E_extra_pc[6]~q ),
	.prn(vcc));
defparam \E_extra_pc[6] .is_wysiwyg = "true";
defparam \E_extra_pc[6] .power_up = "low";

cyclonev_lcell_comb \M_pipe_flush_waddr_nxt[6]~12 (
	.dataa(!\E_src1[8]~19_combout ),
	.datab(!\E_src1[8]~20_combout ),
	.datac(!\E_extra_pc[6]~q ),
	.datad(!\M_pipe_flush_waddr[7]~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_pipe_flush_waddr_nxt[6]~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_pipe_flush_waddr_nxt[6]~12 .extended_lut = "off";
defparam \M_pipe_flush_waddr_nxt[6]~12 .lut_mask = 64'hFAFCFAFCFAFCFAFC;
defparam \M_pipe_flush_waddr_nxt[6]~12 .shared_arith = "off";

cyclonev_lcell_comb \M_pipe_flush_waddr_nxt[6]~13 (
	.dataa(!\E_iw[12]~q ),
	.datab(!\E_hbreak_req~combout ),
	.datac(!\E_ctrl_jmp_indirect~q ),
	.datad(!\E_ctrl_jmp_direct~q ),
	.datae(!\M_pipe_flush_waddr[7]~0_combout ),
	.dataf(!\M_pipe_flush_waddr_nxt[6]~12_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_pipe_flush_waddr_nxt[6]~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_pipe_flush_waddr_nxt[6]~13 .extended_lut = "off";
defparam \M_pipe_flush_waddr_nxt[6]~13 .lut_mask = 64'hFFFFFFFF7FF7FFFF;
defparam \M_pipe_flush_waddr_nxt[6]~13 .shared_arith = "off";

dffeas \D_pc[6] (
	.clk(clk_clk),
	.d(\F_pc[6]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\D_pc[6]~q ),
	.prn(vcc));
defparam \D_pc[6] .is_wysiwyg = "true";
defparam \D_pc[6] .power_up = "low";

dffeas \E_pc[6] (
	.clk(clk_clk),
	.d(\D_pc[6]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_pc[6]~q ),
	.prn(vcc));
defparam \E_pc[6] .is_wysiwyg = "true";
defparam \E_pc[6] .power_up = "low";

dffeas \M_pipe_flush_waddr[6] (
	.clk(clk_clk),
	.d(\M_pipe_flush_waddr_nxt[6]~13_combout ),
	.asdata(\E_pc[6]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\M_pipe_flush_waddr[7]~2_combout ),
	.sload(\E_hbreak_req~combout ),
	.ena(\W_stall~combout ),
	.q(\M_pipe_flush_waddr[6]~q ),
	.prn(vcc));
defparam \M_pipe_flush_waddr[6] .is_wysiwyg = "true";
defparam \M_pipe_flush_waddr[6] .power_up = "low";

cyclonev_lcell_comb \F_ic_tag_rd_addr_nxt[3]~3 (
	.dataa(!\M_pipe_flush_waddr[6]~q ),
	.datab(!\D_pc[6]~q ),
	.datac(!\Add3~45_sumout ),
	.datad(!\D_br_taken_waddr_partial[6]~q ),
	.datae(!\F_ic_data_rd_addr_nxt[0]~0_combout ),
	.dataf(!\F_kill~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ic_tag_rd_addr_nxt[3]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ic_tag_rd_addr_nxt[3]~3 .extended_lut = "off";
defparam \F_ic_tag_rd_addr_nxt[3]~3 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \F_ic_tag_rd_addr_nxt[3]~3 .shared_arith = "off";

dffeas \F_pc[6] (
	.clk(clk_clk),
	.d(\F_ic_tag_rd_addr_nxt[3]~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\F_pc[6]~q ),
	.prn(vcc));
defparam \F_pc[6] .is_wysiwyg = "true";
defparam \F_pc[6] .power_up = "low";

cyclonev_lcell_comb \Add3~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\F_pc[7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~46 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add3~41_sumout ),
	.cout(\Add3~42 ),
	.shareout());
defparam \Add3~41 .extended_lut = "off";
defparam \Add3~41 .lut_mask = 64'h00000000000000FF;
defparam \Add3~41 .shared_arith = "off";

cyclonev_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\processor_cpu_ic_data|the_altsyncram|auto_generated|q_b[15] ),
	.datae(gnd),
	.dataf(!\Add3~41_sumout ),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout());
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~21 .shared_arith = "off";

dffeas \D_br_taken_waddr_partial[7] (
	.clk(clk_clk),
	.d(\Add0~21_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\D_br_taken_waddr_partial[7]~q ),
	.prn(vcc));
defparam \D_br_taken_waddr_partial[7] .is_wysiwyg = "true";
defparam \D_br_taken_waddr_partial[7] .power_up = "low";

dffeas \D_pc_plus_one[7] (
	.clk(clk_clk),
	.d(\Add3~41_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\D_pc_plus_one[7]~q ),
	.prn(vcc));
defparam \D_pc_plus_one[7] .is_wysiwyg = "true";
defparam \D_pc_plus_one[7] .power_up = "low";

dffeas \E_extra_pc[7] (
	.clk(clk_clk),
	.d(\D_br_taken_waddr_partial[7]~q ),
	.asdata(\D_pc_plus_one[7]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\D_br_pred_not_taken~combout ),
	.ena(\W_stall~combout ),
	.q(\E_extra_pc[7]~q ),
	.prn(vcc));
defparam \E_extra_pc[7] .is_wysiwyg = "true";
defparam \E_extra_pc[7] .power_up = "low";

cyclonev_lcell_comb \M_pipe_flush_waddr_nxt[7]~14 (
	.dataa(!\E_src1_hazard_M~q ),
	.datab(!\M_wr_data_unfiltered[9]~6_combout ),
	.datac(!\E_src1_prelim[9]~q ),
	.datad(!\E_extra_pc[7]~q ),
	.datae(!\M_pipe_flush_waddr[7]~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_pipe_flush_waddr_nxt[7]~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_pipe_flush_waddr_nxt[7]~14 .extended_lut = "off";
defparam \M_pipe_flush_waddr_nxt[7]~14 .lut_mask = 64'h7FFFBFFF7FFFBFFF;
defparam \M_pipe_flush_waddr_nxt[7]~14 .shared_arith = "off";

cyclonev_lcell_comb \M_pipe_flush_waddr_nxt[7]~15 (
	.dataa(!\E_iw[13]~q ),
	.datab(!\E_hbreak_req~combout ),
	.datac(!\E_ctrl_jmp_indirect~q ),
	.datad(!\E_ctrl_jmp_direct~q ),
	.datae(!\M_pipe_flush_waddr[7]~0_combout ),
	.dataf(!\M_pipe_flush_waddr_nxt[7]~14_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_pipe_flush_waddr_nxt[7]~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_pipe_flush_waddr_nxt[7]~15 .extended_lut = "off";
defparam \M_pipe_flush_waddr_nxt[7]~15 .lut_mask = 64'h7FF7FFFFFFFFFFFF;
defparam \M_pipe_flush_waddr_nxt[7]~15 .shared_arith = "off";

dffeas \D_pc[7] (
	.clk(clk_clk),
	.d(\F_pc[7]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\D_pc[7]~q ),
	.prn(vcc));
defparam \D_pc[7] .is_wysiwyg = "true";
defparam \D_pc[7] .power_up = "low";

dffeas \E_pc[7] (
	.clk(clk_clk),
	.d(\D_pc[7]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_pc[7]~q ),
	.prn(vcc));
defparam \E_pc[7] .is_wysiwyg = "true";
defparam \E_pc[7] .power_up = "low";

dffeas \M_pipe_flush_waddr[7] (
	.clk(clk_clk),
	.d(\M_pipe_flush_waddr_nxt[7]~15_combout ),
	.asdata(\E_pc[7]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\M_pipe_flush_waddr[7]~2_combout ),
	.sload(\E_hbreak_req~combout ),
	.ena(\W_stall~combout ),
	.q(\M_pipe_flush_waddr[7]~q ),
	.prn(vcc));
defparam \M_pipe_flush_waddr[7] .is_wysiwyg = "true";
defparam \M_pipe_flush_waddr[7] .power_up = "low";

cyclonev_lcell_comb \F_ic_tag_rd_addr_nxt[4]~4 (
	.dataa(!\M_pipe_flush_waddr[7]~q ),
	.datab(!\D_pc[7]~q ),
	.datac(!\Add3~41_sumout ),
	.datad(!\D_br_taken_waddr_partial[7]~q ),
	.datae(!\F_ic_data_rd_addr_nxt[0]~0_combout ),
	.dataf(!\F_kill~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ic_tag_rd_addr_nxt[4]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ic_tag_rd_addr_nxt[4]~4 .extended_lut = "off";
defparam \F_ic_tag_rd_addr_nxt[4]~4 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \F_ic_tag_rd_addr_nxt[4]~4 .shared_arith = "off";

dffeas \F_pc[7] (
	.clk(clk_clk),
	.d(\F_ic_tag_rd_addr_nxt[4]~4_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\F_pc[7]~q ),
	.prn(vcc));
defparam \F_pc[7] .is_wysiwyg = "true";
defparam \F_pc[7] .power_up = "low";

cyclonev_lcell_comb \Add3~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\F_pc[8]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~42 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add3~37_sumout ),
	.cout(\Add3~38 ),
	.shareout());
defparam \Add3~37 .extended_lut = "off";
defparam \Add3~37 .lut_mask = 64'h00000000000000FF;
defparam \Add3~37 .shared_arith = "off";

cyclonev_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\processor_cpu_ic_data|the_altsyncram|auto_generated|q_b[16] ),
	.datae(gnd),
	.dataf(!\Add3~37_sumout ),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout());
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~17 .shared_arith = "off";

dffeas \D_br_taken_waddr_partial[8] (
	.clk(clk_clk),
	.d(\Add0~17_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\D_br_taken_waddr_partial[8]~q ),
	.prn(vcc));
defparam \D_br_taken_waddr_partial[8] .is_wysiwyg = "true";
defparam \D_br_taken_waddr_partial[8] .power_up = "low";

dffeas \D_pc_plus_one[8] (
	.clk(clk_clk),
	.d(\Add3~37_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\D_pc_plus_one[8]~q ),
	.prn(vcc));
defparam \D_pc_plus_one[8] .is_wysiwyg = "true";
defparam \D_pc_plus_one[8] .power_up = "low";

dffeas \E_extra_pc[8] (
	.clk(clk_clk),
	.d(\D_br_taken_waddr_partial[8]~q ),
	.asdata(\D_pc_plus_one[8]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\D_br_pred_not_taken~combout ),
	.ena(\W_stall~combout ),
	.q(\E_extra_pc[8]~q ),
	.prn(vcc));
defparam \E_extra_pc[8] .is_wysiwyg = "true";
defparam \E_extra_pc[8] .power_up = "low";

cyclonev_lcell_comb \M_pipe_flush_waddr_nxt[8]~16 (
	.dataa(!\E_src1[10]~15_combout ),
	.datab(!\E_src1[10]~16_combout ),
	.datac(!\E_extra_pc[8]~q ),
	.datad(!\M_pipe_flush_waddr[7]~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_pipe_flush_waddr_nxt[8]~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_pipe_flush_waddr_nxt[8]~16 .extended_lut = "off";
defparam \M_pipe_flush_waddr_nxt[8]~16 .lut_mask = 64'hFAFCFAFCFAFCFAFC;
defparam \M_pipe_flush_waddr_nxt[8]~16 .shared_arith = "off";

cyclonev_lcell_comb \M_pipe_flush_waddr_nxt[8]~17 (
	.dataa(!\E_iw[14]~q ),
	.datab(!\E_hbreak_req~combout ),
	.datac(!\E_ctrl_jmp_indirect~q ),
	.datad(!\E_ctrl_jmp_direct~q ),
	.datae(!\M_pipe_flush_waddr[7]~0_combout ),
	.dataf(!\M_pipe_flush_waddr_nxt[8]~16_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_pipe_flush_waddr_nxt[8]~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_pipe_flush_waddr_nxt[8]~17 .extended_lut = "off";
defparam \M_pipe_flush_waddr_nxt[8]~17 .lut_mask = 64'hFFFFFFFF7FF7FFFF;
defparam \M_pipe_flush_waddr_nxt[8]~17 .shared_arith = "off";

dffeas \D_pc[8] (
	.clk(clk_clk),
	.d(\F_pc[8]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\D_pc[8]~q ),
	.prn(vcc));
defparam \D_pc[8] .is_wysiwyg = "true";
defparam \D_pc[8] .power_up = "low";

dffeas \E_pc[8] (
	.clk(clk_clk),
	.d(\D_pc[8]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_pc[8]~q ),
	.prn(vcc));
defparam \E_pc[8] .is_wysiwyg = "true";
defparam \E_pc[8] .power_up = "low";

dffeas \M_pipe_flush_waddr[8] (
	.clk(clk_clk),
	.d(\M_pipe_flush_waddr_nxt[8]~17_combout ),
	.asdata(\E_pc[8]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\M_pipe_flush_waddr[7]~2_combout ),
	.sload(\E_hbreak_req~combout ),
	.ena(\W_stall~combout ),
	.q(\M_pipe_flush_waddr[8]~q ),
	.prn(vcc));
defparam \M_pipe_flush_waddr[8] .is_wysiwyg = "true";
defparam \M_pipe_flush_waddr[8] .power_up = "low";

cyclonev_lcell_comb \F_ic_tag_rd_addr_nxt[5]~5 (
	.dataa(!\M_pipe_flush_waddr[8]~q ),
	.datab(!\D_pc[8]~q ),
	.datac(!\Add3~37_sumout ),
	.datad(!\D_br_taken_waddr_partial[8]~q ),
	.datae(!\F_ic_data_rd_addr_nxt[0]~0_combout ),
	.dataf(!\F_kill~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ic_tag_rd_addr_nxt[5]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ic_tag_rd_addr_nxt[5]~5 .extended_lut = "off";
defparam \F_ic_tag_rd_addr_nxt[5]~5 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \F_ic_tag_rd_addr_nxt[5]~5 .shared_arith = "off";

dffeas \F_pc[8] (
	.clk(clk_clk),
	.d(\F_ic_tag_rd_addr_nxt[5]~5_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\F_pc[8]~q ),
	.prn(vcc));
defparam \F_pc[8] .is_wysiwyg = "true";
defparam \F_pc[8] .power_up = "low";

cyclonev_lcell_comb \Add3~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\F_pc[9]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add3~33_sumout ),
	.cout(\Add3~34 ),
	.shareout());
defparam \Add3~33 .extended_lut = "off";
defparam \Add3~33 .lut_mask = 64'h00000000000000FF;
defparam \Add3~33 .shared_arith = "off";

cyclonev_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\processor_cpu_ic_data|the_altsyncram|auto_generated|q_b[17] ),
	.datae(gnd),
	.dataf(!\Add3~33_sumout ),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout());
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~13 .shared_arith = "off";

dffeas \D_br_taken_waddr_partial[9] (
	.clk(clk_clk),
	.d(\Add0~13_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\D_br_taken_waddr_partial[9]~q ),
	.prn(vcc));
defparam \D_br_taken_waddr_partial[9] .is_wysiwyg = "true";
defparam \D_br_taken_waddr_partial[9] .power_up = "low";

dffeas \D_pc_plus_one[9] (
	.clk(clk_clk),
	.d(\Add3~33_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\D_pc_plus_one[9]~q ),
	.prn(vcc));
defparam \D_pc_plus_one[9] .is_wysiwyg = "true";
defparam \D_pc_plus_one[9] .power_up = "low";

dffeas \E_extra_pc[9] (
	.clk(clk_clk),
	.d(\D_br_taken_waddr_partial[9]~q ),
	.asdata(\D_pc_plus_one[9]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\D_br_pred_not_taken~combout ),
	.ena(\W_stall~combout ),
	.q(\E_extra_pc[9]~q ),
	.prn(vcc));
defparam \E_extra_pc[9] .is_wysiwyg = "true";
defparam \E_extra_pc[9] .power_up = "low";

cyclonev_lcell_comb \M_pipe_flush_waddr[7]~3 (
	.dataa(!\E_hbreak_req~combout ),
	.datab(!\E_ctrl_jmp_indirect~q ),
	.datac(!\E_ctrl_jmp_direct~q ),
	.datad(!\M_pipe_flush_waddr[7]~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_pipe_flush_waddr[7]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_pipe_flush_waddr[7]~3 .extended_lut = "off";
defparam \M_pipe_flush_waddr[7]~3 .lut_mask = 64'hFFEFFFEFFFEFFFEF;
defparam \M_pipe_flush_waddr[7]~3 .shared_arith = "off";

cyclonev_lcell_comb \M_pipe_flush_waddr_nxt[9]~23 (
	.dataa(!\E_extra_pc[9]~q ),
	.datab(!\E_src1[11]~14_combout ),
	.datac(!\E_ctrl_exception~q ),
	.datad(!\E_iw[15]~q ),
	.datae(!\M_pipe_flush_waddr[7]~1_combout ),
	.dataf(!\M_pipe_flush_waddr[7]~3_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_pipe_flush_waddr_nxt[9]~23_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_pipe_flush_waddr_nxt[9]~23 .extended_lut = "off";
defparam \M_pipe_flush_waddr_nxt[9]~23 .lut_mask = 64'hF7FFFFFFFFFFF7FF;
defparam \M_pipe_flush_waddr_nxt[9]~23 .shared_arith = "off";

dffeas \D_pc[9] (
	.clk(clk_clk),
	.d(\F_pc[9]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\D_pc[9]~q ),
	.prn(vcc));
defparam \D_pc[9] .is_wysiwyg = "true";
defparam \D_pc[9] .power_up = "low";

dffeas \E_pc[9] (
	.clk(clk_clk),
	.d(\D_pc[9]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_pc[9]~q ),
	.prn(vcc));
defparam \E_pc[9] .is_wysiwyg = "true";
defparam \E_pc[9] .power_up = "low";

dffeas \M_pipe_flush_waddr[9] (
	.clk(clk_clk),
	.d(\M_pipe_flush_waddr_nxt[9]~23_combout ),
	.asdata(\E_pc[9]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\M_pipe_flush_waddr[7]~2_combout ),
	.sload(\E_hbreak_req~combout ),
	.ena(\W_stall~combout ),
	.q(\M_pipe_flush_waddr[9]~q ),
	.prn(vcc));
defparam \M_pipe_flush_waddr[9] .is_wysiwyg = "true";
defparam \M_pipe_flush_waddr[9] .power_up = "low";

cyclonev_lcell_comb \F_pc_nxt[9]~3 (
	.dataa(!\M_pipe_flush_waddr[9]~q ),
	.datab(!\D_pc[9]~q ),
	.datac(!\Add3~33_sumout ),
	.datad(!\D_br_taken_waddr_partial[9]~q ),
	.datae(!\F_ic_data_rd_addr_nxt[0]~0_combout ),
	.dataf(!\F_kill~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_pc_nxt[9]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_pc_nxt[9]~3 .extended_lut = "off";
defparam \F_pc_nxt[9]~3 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \F_pc_nxt[9]~3 .shared_arith = "off";

dffeas \F_pc[9] (
	.clk(clk_clk),
	.d(\F_pc_nxt[9]~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\F_pc[9]~q ),
	.prn(vcc));
defparam \F_pc[9] .is_wysiwyg = "true";
defparam \F_pc[9] .power_up = "low";

cyclonev_lcell_comb \Add3~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\F_pc[10]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add3~29_sumout ),
	.cout(\Add3~30 ),
	.shareout());
defparam \Add3~29 .extended_lut = "off";
defparam \Add3~29 .lut_mask = 64'h00000000000000FF;
defparam \Add3~29 .shared_arith = "off";

dffeas \D_pc_plus_one[10] (
	.clk(clk_clk),
	.d(\Add3~29_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\D_pc_plus_one[10]~q ),
	.prn(vcc));
defparam \D_pc_plus_one[10] .is_wysiwyg = "true";
defparam \D_pc_plus_one[10] .power_up = "low";

cyclonev_lcell_comb \Add0~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~41_sumout ),
	.cout(),
	.shareout());
defparam \Add0~41 .extended_lut = "off";
defparam \Add0~41 .lut_mask = 64'h0000000000000000;
defparam \Add0~41 .shared_arith = "off";

dffeas \D_br_taken_waddr_partial[10] (
	.clk(clk_clk),
	.d(\Add0~41_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\D_br_taken_waddr_partial[10]~q ),
	.prn(vcc));
defparam \D_br_taken_waddr_partial[10] .is_wysiwyg = "true";
defparam \D_br_taken_waddr_partial[10] .power_up = "low";

cyclonev_lcell_comb \Add1~22 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\D_br_taken_waddr_partial[10]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\Add1~22_cout ),
	.shareout());
defparam \Add1~22 .extended_lut = "off";
defparam \Add1~22 .lut_mask = 64'h00000000000000FF;
defparam \Add1~22 .shared_arith = "off";

cyclonev_lcell_comb \Add1~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\D_pc_plus_one[10]~q ),
	.datae(gnd),
	.dataf(!\D_iw[18]~q ),
	.datag(gnd),
	.cin(\Add1~22_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~17_sumout ),
	.cout(\Add1~18 ),
	.shareout());
defparam \Add1~17 .extended_lut = "off";
defparam \Add1~17 .lut_mask = 64'h0000FF00000000FF;
defparam \Add1~17 .shared_arith = "off";

dffeas \E_extra_pc[10] (
	.clk(clk_clk),
	.d(\Add1~17_sumout ),
	.asdata(\D_pc_plus_one[10]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\D_br_pred_not_taken~combout ),
	.ena(\W_stall~combout ),
	.q(\E_extra_pc[10]~q ),
	.prn(vcc));
defparam \E_extra_pc[10] .is_wysiwyg = "true";
defparam \E_extra_pc[10] .power_up = "low";

cyclonev_lcell_comb \M_pipe_flush_waddr_nxt[10]~19 (
	.dataa(!\E_src1_hazard_M~q ),
	.datab(!\E_extra_pc[10]~q ),
	.datac(!\M_wr_data_unfiltered[12]~4_combout ),
	.datad(!\E_src1_prelim[12]~q ),
	.datae(!\M_pipe_flush_waddr[7]~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_pipe_flush_waddr_nxt[10]~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_pipe_flush_waddr_nxt[10]~19 .extended_lut = "off";
defparam \M_pipe_flush_waddr_nxt[10]~19 .lut_mask = 64'h7FFFBFFF7FFFBFFF;
defparam \M_pipe_flush_waddr_nxt[10]~19 .shared_arith = "off";

cyclonev_lcell_comb \M_pipe_flush_waddr_nxt[10]~20 (
	.dataa(!\E_iw[16]~q ),
	.datab(!\E_hbreak_req~combout ),
	.datac(!\E_ctrl_jmp_indirect~q ),
	.datad(!\E_ctrl_jmp_direct~q ),
	.datae(!\M_pipe_flush_waddr[7]~0_combout ),
	.dataf(!\M_pipe_flush_waddr_nxt[10]~19_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_pipe_flush_waddr_nxt[10]~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_pipe_flush_waddr_nxt[10]~20 .extended_lut = "off";
defparam \M_pipe_flush_waddr_nxt[10]~20 .lut_mask = 64'h7FF7FFFFFFFFFFFF;
defparam \M_pipe_flush_waddr_nxt[10]~20 .shared_arith = "off";

dffeas \D_pc[10] (
	.clk(clk_clk),
	.d(\F_pc[10]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\D_pc[10]~q ),
	.prn(vcc));
defparam \D_pc[10] .is_wysiwyg = "true";
defparam \D_pc[10] .power_up = "low";

dffeas \E_pc[10] (
	.clk(clk_clk),
	.d(\D_pc[10]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_pc[10]~q ),
	.prn(vcc));
defparam \E_pc[10] .is_wysiwyg = "true";
defparam \E_pc[10] .power_up = "low";

dffeas \M_pipe_flush_waddr[10] (
	.clk(clk_clk),
	.d(\M_pipe_flush_waddr_nxt[10]~20_combout ),
	.asdata(\E_pc[10]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\M_pipe_flush_waddr[7]~2_combout ),
	.sload(\E_hbreak_req~combout ),
	.ena(\W_stall~combout ),
	.q(\M_pipe_flush_waddr[10]~q ),
	.prn(vcc));
defparam \M_pipe_flush_waddr[10] .is_wysiwyg = "true";
defparam \M_pipe_flush_waddr[10] .power_up = "low";

cyclonev_lcell_comb \F_pc_nxt[10]~1 (
	.dataa(!\M_pipe_flush_waddr[10]~q ),
	.datab(!\D_pc[10]~q ),
	.datac(!\Add3~29_sumout ),
	.datad(!\Add1~17_sumout ),
	.datae(!\F_ic_data_rd_addr_nxt[0]~0_combout ),
	.dataf(!\F_kill~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_pc_nxt[10]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_pc_nxt[10]~1 .extended_lut = "off";
defparam \F_pc_nxt[10]~1 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \F_pc_nxt[10]~1 .shared_arith = "off";

dffeas \F_pc[10] (
	.clk(clk_clk),
	.d(\F_pc_nxt[10]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\F_pc[10]~q ),
	.prn(vcc));
defparam \F_pc[10] .is_wysiwyg = "true";
defparam \F_pc[10] .power_up = "low";

cyclonev_lcell_comb \Add3~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\F_pc[11]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add3~25_sumout ),
	.cout(\Add3~26 ),
	.shareout());
defparam \Add3~25 .extended_lut = "off";
defparam \Add3~25 .lut_mask = 64'h00000000000000FF;
defparam \Add3~25 .shared_arith = "off";

dffeas \D_pc_plus_one[11] (
	.clk(clk_clk),
	.d(\Add3~25_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\D_pc_plus_one[11]~q ),
	.prn(vcc));
defparam \D_pc_plus_one[11] .is_wysiwyg = "true";
defparam \D_pc_plus_one[11] .power_up = "low";

cyclonev_lcell_comb \Add1~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\D_pc_plus_one[11]~q ),
	.datae(gnd),
	.dataf(!\D_iw[19]~q ),
	.datag(gnd),
	.cin(\Add1~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~13_sumout ),
	.cout(\Add1~14 ),
	.shareout());
defparam \Add1~13 .extended_lut = "off";
defparam \Add1~13 .lut_mask = 64'h0000FF00000000FF;
defparam \Add1~13 .shared_arith = "off";

dffeas \E_extra_pc[11] (
	.clk(clk_clk),
	.d(\Add1~13_sumout ),
	.asdata(\D_pc_plus_one[11]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\D_br_pred_not_taken~combout ),
	.ena(\W_stall~combout ),
	.q(\E_extra_pc[11]~q ),
	.prn(vcc));
defparam \E_extra_pc[11] .is_wysiwyg = "true";
defparam \E_extra_pc[11] .power_up = "low";

cyclonev_lcell_comb \M_pipe_flush_waddr_nxt[11]~24 (
	.dataa(!\E_src1_hazard_M~q ),
	.datab(!\M_wr_data_unfiltered[13]~3_combout ),
	.datac(!\E_src1_prelim[13]~q ),
	.datad(!\E_extra_pc[11]~q ),
	.datae(!\M_pipe_flush_waddr[7]~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_pipe_flush_waddr_nxt[11]~24_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_pipe_flush_waddr_nxt[11]~24 .extended_lut = "off";
defparam \M_pipe_flush_waddr_nxt[11]~24 .lut_mask = 64'h7FFFBFFF7FFFBFFF;
defparam \M_pipe_flush_waddr_nxt[11]~24 .shared_arith = "off";

dffeas \E_iw[17] (
	.clk(clk_clk),
	.d(\D_iw[17]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_iw[17]~q ),
	.prn(vcc));
defparam \E_iw[17] .is_wysiwyg = "true";
defparam \E_iw[17] .power_up = "low";

cyclonev_lcell_comb \M_pipe_flush_waddr_nxt[11]~25 (
	.dataa(!\E_hbreak_req~combout ),
	.datab(!\E_ctrl_jmp_indirect~q ),
	.datac(!\E_ctrl_jmp_direct~q ),
	.datad(!\M_pipe_flush_waddr[7]~0_combout ),
	.datae(!\M_pipe_flush_waddr_nxt[11]~24_combout ),
	.dataf(!\E_iw[17]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_pipe_flush_waddr_nxt[11]~25_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_pipe_flush_waddr_nxt[11]~25 .extended_lut = "off";
defparam \M_pipe_flush_waddr_nxt[11]~25 .lut_mask = 64'h7DFFFFFFFFFFFFFF;
defparam \M_pipe_flush_waddr_nxt[11]~25 .shared_arith = "off";

dffeas \D_pc[11] (
	.clk(clk_clk),
	.d(\F_pc[11]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\D_pc[11]~q ),
	.prn(vcc));
defparam \D_pc[11] .is_wysiwyg = "true";
defparam \D_pc[11] .power_up = "low";

dffeas \E_pc[11] (
	.clk(clk_clk),
	.d(\D_pc[11]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_pc[11]~q ),
	.prn(vcc));
defparam \E_pc[11] .is_wysiwyg = "true";
defparam \E_pc[11] .power_up = "low";

dffeas \M_pipe_flush_waddr[11] (
	.clk(clk_clk),
	.d(\M_pipe_flush_waddr_nxt[11]~25_combout ),
	.asdata(\E_pc[11]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\M_pipe_flush_waddr[7]~2_combout ),
	.sload(\E_hbreak_req~combout ),
	.ena(\W_stall~combout ),
	.q(\M_pipe_flush_waddr[11]~q ),
	.prn(vcc));
defparam \M_pipe_flush_waddr[11] .is_wysiwyg = "true";
defparam \M_pipe_flush_waddr[11] .power_up = "low";

cyclonev_lcell_comb \F_pc_nxt[11]~4 (
	.dataa(!\M_pipe_flush_waddr[11]~q ),
	.datab(!\D_pc[11]~q ),
	.datac(!\Add3~25_sumout ),
	.datad(!\Add1~13_sumout ),
	.datae(!\F_ic_data_rd_addr_nxt[0]~0_combout ),
	.dataf(!\F_kill~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_pc_nxt[11]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_pc_nxt[11]~4 .extended_lut = "off";
defparam \F_pc_nxt[11]~4 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \F_pc_nxt[11]~4 .shared_arith = "off";

dffeas \F_pc[11] (
	.clk(clk_clk),
	.d(\F_pc_nxt[11]~4_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\F_pc[11]~q ),
	.prn(vcc));
defparam \F_pc[11] .is_wysiwyg = "true";
defparam \F_pc[11] .power_up = "low";

cyclonev_lcell_comb \Add3~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\F_pc[12]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add3~21_sumout ),
	.cout(\Add3~22 ),
	.shareout());
defparam \Add3~21 .extended_lut = "off";
defparam \Add3~21 .lut_mask = 64'h00000000000000FF;
defparam \Add3~21 .shared_arith = "off";

dffeas \D_pc_plus_one[12] (
	.clk(clk_clk),
	.d(\Add3~21_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\D_pc_plus_one[12]~q ),
	.prn(vcc));
defparam \D_pc_plus_one[12] .is_wysiwyg = "true";
defparam \D_pc_plus_one[12] .power_up = "low";

cyclonev_lcell_comb \Add1~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\D_pc_plus_one[12]~q ),
	.datae(gnd),
	.dataf(!\D_iw[20]~q ),
	.datag(gnd),
	.cin(\Add1~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~9_sumout ),
	.cout(\Add1~10 ),
	.shareout());
defparam \Add1~9 .extended_lut = "off";
defparam \Add1~9 .lut_mask = 64'h0000FF00000000FF;
defparam \Add1~9 .shared_arith = "off";

dffeas \E_extra_pc[12] (
	.clk(clk_clk),
	.d(\Add1~9_sumout ),
	.asdata(\D_pc_plus_one[12]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\D_br_pred_not_taken~combout ),
	.ena(\W_stall~combout ),
	.q(\E_extra_pc[12]~q ),
	.prn(vcc));
defparam \E_extra_pc[12] .is_wysiwyg = "true";
defparam \E_extra_pc[12] .power_up = "low";

cyclonev_lcell_comb \M_pipe_flush_waddr_nxt[12]~26 (
	.dataa(!\E_src1_hazard_M~q ),
	.datab(!\M_wr_data_unfiltered[14]~2_combout ),
	.datac(!\E_src1_prelim[14]~q ),
	.datad(!\E_extra_pc[12]~q ),
	.datae(!\M_pipe_flush_waddr[7]~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_pipe_flush_waddr_nxt[12]~26_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_pipe_flush_waddr_nxt[12]~26 .extended_lut = "off";
defparam \M_pipe_flush_waddr_nxt[12]~26 .lut_mask = 64'h7FFFBFFF7FFFBFFF;
defparam \M_pipe_flush_waddr_nxt[12]~26 .shared_arith = "off";

dffeas \E_iw[18] (
	.clk(clk_clk),
	.d(\D_iw[18]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_iw[18]~q ),
	.prn(vcc));
defparam \E_iw[18] .is_wysiwyg = "true";
defparam \E_iw[18] .power_up = "low";

cyclonev_lcell_comb \M_pipe_flush_waddr_nxt[12]~27 (
	.dataa(!\E_hbreak_req~combout ),
	.datab(!\E_ctrl_jmp_indirect~q ),
	.datac(!\E_ctrl_jmp_direct~q ),
	.datad(!\M_pipe_flush_waddr[7]~0_combout ),
	.datae(!\M_pipe_flush_waddr_nxt[12]~26_combout ),
	.dataf(!\E_iw[18]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_pipe_flush_waddr_nxt[12]~27_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_pipe_flush_waddr_nxt[12]~27 .extended_lut = "off";
defparam \M_pipe_flush_waddr_nxt[12]~27 .lut_mask = 64'h7DFFFFFFFFFFFFFF;
defparam \M_pipe_flush_waddr_nxt[12]~27 .shared_arith = "off";

dffeas \D_pc[12] (
	.clk(clk_clk),
	.d(\F_pc[12]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\D_pc[12]~q ),
	.prn(vcc));
defparam \D_pc[12] .is_wysiwyg = "true";
defparam \D_pc[12] .power_up = "low";

dffeas \E_pc[12] (
	.clk(clk_clk),
	.d(\D_pc[12]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_pc[12]~q ),
	.prn(vcc));
defparam \E_pc[12] .is_wysiwyg = "true";
defparam \E_pc[12] .power_up = "low";

dffeas \M_pipe_flush_waddr[12] (
	.clk(clk_clk),
	.d(\M_pipe_flush_waddr_nxt[12]~27_combout ),
	.asdata(\E_pc[12]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\M_pipe_flush_waddr[7]~2_combout ),
	.sload(\E_hbreak_req~combout ),
	.ena(\W_stall~combout ),
	.q(\M_pipe_flush_waddr[12]~q ),
	.prn(vcc));
defparam \M_pipe_flush_waddr[12] .is_wysiwyg = "true";
defparam \M_pipe_flush_waddr[12] .power_up = "low";

cyclonev_lcell_comb \F_pc_nxt[12]~5 (
	.dataa(!\M_pipe_flush_waddr[12]~q ),
	.datab(!\D_pc[12]~q ),
	.datac(!\Add3~21_sumout ),
	.datad(!\Add1~9_sumout ),
	.datae(!\F_ic_data_rd_addr_nxt[0]~0_combout ),
	.dataf(!\F_kill~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_pc_nxt[12]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_pc_nxt[12]~5 .extended_lut = "off";
defparam \F_pc_nxt[12]~5 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \F_pc_nxt[12]~5 .shared_arith = "off";

dffeas \F_pc[12] (
	.clk(clk_clk),
	.d(\F_pc_nxt[12]~5_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\F_pc[12]~q ),
	.prn(vcc));
defparam \F_pc[12] .is_wysiwyg = "true";
defparam \F_pc[12] .power_up = "low";

cyclonev_lcell_comb \Add3~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\F_pc[13]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add3~17_sumout ),
	.cout(\Add3~18 ),
	.shareout());
defparam \Add3~17 .extended_lut = "off";
defparam \Add3~17 .lut_mask = 64'h00000000000000FF;
defparam \Add3~17 .shared_arith = "off";

dffeas \D_pc_plus_one[13] (
	.clk(clk_clk),
	.d(\Add3~17_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\D_pc_plus_one[13]~q ),
	.prn(vcc));
defparam \D_pc_plus_one[13] .is_wysiwyg = "true";
defparam \D_pc_plus_one[13] .power_up = "low";

cyclonev_lcell_comb \Add1~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\D_pc_plus_one[13]~q ),
	.datae(gnd),
	.dataf(!\D_iw[21]~q ),
	.datag(gnd),
	.cin(\Add1~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~5_sumout ),
	.cout(\Add1~6 ),
	.shareout());
defparam \Add1~5 .extended_lut = "off";
defparam \Add1~5 .lut_mask = 64'h0000FF00000000FF;
defparam \Add1~5 .shared_arith = "off";

dffeas \E_extra_pc[13] (
	.clk(clk_clk),
	.d(\Add1~5_sumout ),
	.asdata(\D_pc_plus_one[13]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\D_br_pred_not_taken~combout ),
	.ena(\W_stall~combout ),
	.q(\E_extra_pc[13]~q ),
	.prn(vcc));
defparam \E_extra_pc[13] .is_wysiwyg = "true";
defparam \E_extra_pc[13] .power_up = "low";

dffeas \E_iw[19] (
	.clk(clk_clk),
	.d(\D_iw[19]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_iw[19]~q ),
	.prn(vcc));
defparam \E_iw[19] .is_wysiwyg = "true";
defparam \E_iw[19] .power_up = "low";

cyclonev_lcell_comb \M_pipe_flush_waddr_nxt[13]~21 (
	.dataa(!\E_extra_pc[13]~q ),
	.datab(!\E_ctrl_break~q ),
	.datac(!\E_ctrl_exception~q ),
	.datad(!\E_ctrl_crst~q ),
	.datae(!\E_ctrl_jmp_direct~q ),
	.dataf(!\E_iw[19]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_pipe_flush_waddr_nxt[13]~21_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_pipe_flush_waddr_nxt[13]~21 .extended_lut = "off";
defparam \M_pipe_flush_waddr_nxt[13]~21 .lut_mask = 64'hFFFFFFFFFFBBFFF3;
defparam \M_pipe_flush_waddr_nxt[13]~21 .shared_arith = "off";

cyclonev_lcell_comb \M_pipe_flush_waddr_nxt[13]~22 (
	.dataa(!\E_hbreak_req~combout ),
	.datab(!\E_src1[15]~10_combout ),
	.datac(!\E_ctrl_jmp_indirect~q ),
	.datad(!\E_pc[13]~q ),
	.datae(!\M_pipe_flush_waddr_nxt[13]~21_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_pipe_flush_waddr_nxt[13]~22_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_pipe_flush_waddr_nxt[13]~22 .extended_lut = "off";
defparam \M_pipe_flush_waddr_nxt[13]~22 .lut_mask = 64'hFFDEFFFFFFDEFFFF;
defparam \M_pipe_flush_waddr_nxt[13]~22 .shared_arith = "off";

dffeas \M_pipe_flush_waddr[13] (
	.clk(clk_clk),
	.d(\M_pipe_flush_waddr_nxt[13]~22_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\M_pipe_flush_waddr[13]~q ),
	.prn(vcc));
defparam \M_pipe_flush_waddr[13] .is_wysiwyg = "true";
defparam \M_pipe_flush_waddr[13] .power_up = "low";

cyclonev_lcell_comb \F_pc_nxt[13]~2 (
	.dataa(!\M_pipe_flush_waddr[13]~q ),
	.datab(!\D_pc[13]~q ),
	.datac(!\Add3~17_sumout ),
	.datad(!\Add1~5_sumout ),
	.datae(!\F_ic_data_rd_addr_nxt[0]~0_combout ),
	.dataf(!\F_kill~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_pc_nxt[13]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_pc_nxt[13]~2 .extended_lut = "off";
defparam \F_pc_nxt[13]~2 .lut_mask = 64'hBFFFFFFFFFFFBFFF;
defparam \F_pc_nxt[13]~2 .shared_arith = "off";

dffeas \F_pc[13] (
	.clk(clk_clk),
	.d(\F_pc_nxt[13]~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\F_pc[13]~q ),
	.prn(vcc));
defparam \F_pc[13] .is_wysiwyg = "true";
defparam \F_pc[13] .power_up = "low";

cyclonev_lcell_comb \Add3~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\F_pc[14]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add3~13_sumout ),
	.cout(),
	.shareout());
defparam \Add3~13 .extended_lut = "off";
defparam \Add3~13 .lut_mask = 64'h00000000000000FF;
defparam \Add3~13 .shared_arith = "off";

dffeas \D_pc_plus_one[14] (
	.clk(clk_clk),
	.d(\Add3~13_sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\D_pc_plus_one[14]~q ),
	.prn(vcc));
defparam \D_pc_plus_one[14] .is_wysiwyg = "true";
defparam \D_pc_plus_one[14] .power_up = "low";

cyclonev_lcell_comb \Add1~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\D_pc_plus_one[14]~q ),
	.datae(gnd),
	.dataf(!\D_iw[21]~q ),
	.datag(gnd),
	.cin(\Add1~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~1_sumout ),
	.cout(),
	.shareout());
defparam \Add1~1 .extended_lut = "off";
defparam \Add1~1 .lut_mask = 64'h0000FF00000000FF;
defparam \Add1~1 .shared_arith = "off";

dffeas \E_extra_pc[14] (
	.clk(clk_clk),
	.d(\Add1~1_sumout ),
	.asdata(\D_pc_plus_one[14]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(\D_br_pred_not_taken~combout ),
	.ena(\W_stall~combout ),
	.q(\E_extra_pc[14]~q ),
	.prn(vcc));
defparam \E_extra_pc[14] .is_wysiwyg = "true";
defparam \E_extra_pc[14] .power_up = "low";

dffeas \E_iw[20] (
	.clk(clk_clk),
	.d(\D_iw[20]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_iw[20]~q ),
	.prn(vcc));
defparam \E_iw[20] .is_wysiwyg = "true";
defparam \E_iw[20] .power_up = "low";

cyclonev_lcell_comb \M_pipe_flush_waddr_nxt[14]~18 (
	.dataa(!\E_extra_pc[14]~q ),
	.datab(!\E_src1[16]~9_combout ),
	.datac(!\E_ctrl_exception~q ),
	.datad(!\E_iw[20]~q ),
	.datae(!\M_pipe_flush_waddr[7]~1_combout ),
	.dataf(!\M_pipe_flush_waddr[7]~3_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_pipe_flush_waddr_nxt[14]~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_pipe_flush_waddr_nxt[14]~18 .extended_lut = "off";
defparam \M_pipe_flush_waddr_nxt[14]~18 .lut_mask = 64'hF7FFFFFFFFFFF7FF;
defparam \M_pipe_flush_waddr_nxt[14]~18 .shared_arith = "off";

dffeas \D_pc[14] (
	.clk(clk_clk),
	.d(\F_pc[14]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\D_pc[14]~q ),
	.prn(vcc));
defparam \D_pc[14] .is_wysiwyg = "true";
defparam \D_pc[14] .power_up = "low";

dffeas \E_pc[14] (
	.clk(clk_clk),
	.d(\D_pc[14]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_pc[14]~q ),
	.prn(vcc));
defparam \E_pc[14] .is_wysiwyg = "true";
defparam \E_pc[14] .power_up = "low";

dffeas \M_pipe_flush_waddr[14] (
	.clk(clk_clk),
	.d(\M_pipe_flush_waddr_nxt[14]~18_combout ),
	.asdata(\E_pc[14]~q ),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\M_pipe_flush_waddr[7]~2_combout ),
	.sload(\E_hbreak_req~combout ),
	.ena(\W_stall~combout ),
	.q(\M_pipe_flush_waddr[14]~q ),
	.prn(vcc));
defparam \M_pipe_flush_waddr[14] .is_wysiwyg = "true";
defparam \M_pipe_flush_waddr[14] .power_up = "low";

cyclonev_lcell_comb \F_pc_nxt[14]~0 (
	.dataa(!\M_pipe_flush_waddr[14]~q ),
	.datab(!\D_pc[14]~q ),
	.datac(!\Add3~13_sumout ),
	.datad(!\Add1~1_sumout ),
	.datae(!\F_ic_data_rd_addr_nxt[0]~0_combout ),
	.dataf(!\F_kill~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_pc_nxt[14]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_pc_nxt[14]~0 .extended_lut = "off";
defparam \F_pc_nxt[14]~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \F_pc_nxt[14]~0 .shared_arith = "off";

dffeas \F_pc[14] (
	.clk(clk_clk),
	.d(\F_pc_nxt[14]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\F_pc[14]~q ),
	.prn(vcc));
defparam \F_pc[14] .is_wysiwyg = "true";
defparam \F_pc[14] .power_up = "low";

cyclonev_lcell_comb \W_valid~0 (
	.dataa(!\M_valid_from_E~q ),
	.datab(!d_write1),
	.datac(!d_read1),
	.datad(!WideOr1),
	.datae(!read_accepted),
	.dataf(!\W_stall~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\W_valid~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \W_valid~0 .extended_lut = "off";
defparam \W_valid~0 .lut_mask = 64'hDFD5FFFFFFFFFFFF;
defparam \W_valid~0 .shared_arith = "off";

dffeas W_valid(
	.clk(clk_clk),
	.d(\W_valid~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_valid~q ),
	.prn(vcc));
defparam W_valid.is_wysiwyg = "true";
defparam W_valid.power_up = "low";

dffeas M_ctrl_crst(
	.clk(clk_clk),
	.d(\E_ctrl_crst~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\M_ctrl_crst~q ),
	.prn(vcc));
defparam M_ctrl_crst.is_wysiwyg = "true";
defparam M_ctrl_crst.power_up = "low";

dffeas W_ctrl_crst(
	.clk(clk_clk),
	.d(\M_ctrl_crst~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\W_ctrl_crst~q ),
	.prn(vcc));
defparam W_ctrl_crst.is_wysiwyg = "true";
defparam W_ctrl_crst.power_up = "low";

cyclonev_lcell_comb \F_inst_ram_hit~0 (
	.dataa(!\W_valid~q ),
	.datab(!\W_ctrl_crst~q ),
	.datac(!\F_pc[9]~q ),
	.datad(!\processor_cpu_ic_tag|the_altsyncram|auto_generated|q_b[0] ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_inst_ram_hit~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_inst_ram_hit~0 .extended_lut = "off";
defparam \F_inst_ram_hit~0 .lut_mask = 64'hEFFEEFFEEFFEEFFE;
defparam \F_inst_ram_hit~0 .shared_arith = "off";

cyclonev_lcell_comb \F_inst_ram_hit~1 (
	.dataa(!\F_pc[11]~q ),
	.datab(!\processor_cpu_ic_tag|the_altsyncram|auto_generated|q_b[2] ),
	.datac(!\F_pc[12]~q ),
	.datad(!\processor_cpu_ic_tag|the_altsyncram|auto_generated|q_b[3] ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_inst_ram_hit~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_inst_ram_hit~1 .extended_lut = "off";
defparam \F_inst_ram_hit~1 .lut_mask = 64'h6996699669966996;
defparam \F_inst_ram_hit~1 .shared_arith = "off";

cyclonev_lcell_comb \F_inst_ram_hit~2 (
	.dataa(!\F_pc[10]~q ),
	.datab(!\processor_cpu_ic_tag|the_altsyncram|auto_generated|q_b[1] ),
	.datac(!\F_pc[13]~q ),
	.datad(!\processor_cpu_ic_tag|the_altsyncram|auto_generated|q_b[4] ),
	.datae(!\F_inst_ram_hit~0_combout ),
	.dataf(!\F_inst_ram_hit~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_inst_ram_hit~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_inst_ram_hit~2 .extended_lut = "off";
defparam \F_inst_ram_hit~2 .lut_mask = 64'h6996FFFFFFFFFFFF;
defparam \F_inst_ram_hit~2 .shared_arith = "off";

cyclonev_lcell_comb \F_inst_ram_hit~3 (
	.dataa(!\F_ic_valid~0_combout ),
	.datab(!\F_pc[14]~q ),
	.datac(!\processor_cpu_ic_tag|the_altsyncram|auto_generated|q_b[5] ),
	.datad(!\F_inst_ram_hit~2_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_inst_ram_hit~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_inst_ram_hit~3 .extended_lut = "off";
defparam \F_inst_ram_hit~3 .lut_mask = 64'h7DFF7DFF7DFF7DFF;
defparam \F_inst_ram_hit~3 .shared_arith = "off";

dffeas D_iw_valid(
	.clk(clk_clk),
	.d(\F_inst_ram_hit~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\D_iw_valid~q ),
	.prn(vcc));
defparam D_iw_valid.is_wysiwyg = "true";
defparam D_iw_valid.power_up = "low";

dffeas D_kill(
	.clk(clk_clk),
	.d(\F_kill~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\D_kill~q ),
	.prn(vcc));
defparam D_kill.is_wysiwyg = "true";
defparam D_kill.power_up = "low";

cyclonev_lcell_comb \D_refetch~0 (
	.dataa(!\D_iw_valid~q ),
	.datab(!\D_kill~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_refetch~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_refetch~0 .extended_lut = "off";
defparam \D_refetch~0 .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \D_refetch~0 .shared_arith = "off";

cyclonev_lcell_comb \F_kill~0 (
	.dataa(!\M_pipe_flush~q ),
	.datab(!\D_refetch~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_kill~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_kill~0 .extended_lut = "off";
defparam \F_kill~0 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \F_kill~0 .shared_arith = "off";

cyclonev_lcell_comb \F_kill~1 (
	.dataa(!\D_iw[21]~q ),
	.datab(!\D_valid~combout ),
	.datac(!\D_ctrl_br~0_combout ),
	.datad(!\Equal4~12_combout ),
	.datae(!\F_kill~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_kill~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_kill~1 .extended_lut = "off";
defparam \F_kill~1 .lut_mask = 64'hFFFF7FFFFFFF7FFF;
defparam \F_kill~1 .shared_arith = "off";

cyclonev_lcell_comb F_issue(
	.dataa(!\F_kill~1_combout ),
	.datab(!\F_ic_valid~0_combout ),
	.datac(!\F_pc[14]~q ),
	.datad(!\processor_cpu_ic_tag|the_altsyncram|auto_generated|q_b[5] ),
	.datae(!\F_inst_ram_hit~2_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_issue~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam F_issue.extended_lut = "off";
defparam F_issue.lut_mask = 64'hBFFBFFFFBFFBFFFF;
defparam F_issue.shared_arith = "off";

dffeas D_issue(
	.clk(clk_clk),
	.d(\F_issue~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\D_issue~q ),
	.prn(vcc));
defparam D_issue.is_wysiwyg = "true";
defparam D_issue.power_up = "low";

cyclonev_lcell_comb D_valid(
	.dataa(!\M_pipe_flush~q ),
	.datab(!\D_issue~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_valid~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam D_valid.extended_lut = "off";
defparam D_valid.lut_mask = 64'h7777777777777777;
defparam D_valid.shared_arith = "off";

dffeas E_valid_from_D(
	.clk(clk_clk),
	.d(\D_valid~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_valid_from_D~q ),
	.prn(vcc));
defparam E_valid_from_D.is_wysiwyg = "true";
defparam E_valid_from_D.power_up = "low";

cyclonev_lcell_comb \E_valid~0 (
	.dataa(!\E_valid_from_D~q ),
	.datab(!\M_pipe_flush~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_valid~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_valid~0 .extended_lut = "off";
defparam \E_valid~0 .lut_mask = 64'h7777777777777777;
defparam \E_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \latched_oci_tb_hbreak_req_next~0 (
	.dataa(!\E_valid~0_combout ),
	.datab(!hbreak_enabled1),
	.datac(!\latched_oci_tb_hbreak_req~q ),
	.datad(!\hbreak_req~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\latched_oci_tb_hbreak_req_next~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \latched_oci_tb_hbreak_req_next~0 .extended_lut = "off";
defparam \latched_oci_tb_hbreak_req_next~0 .lut_mask = 64'hC5FFC5FFC5FFC5FF;
defparam \latched_oci_tb_hbreak_req_next~0 .shared_arith = "off";

dffeas latched_oci_tb_hbreak_req(
	.clk(clk_clk),
	.d(\latched_oci_tb_hbreak_req_next~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\latched_oci_tb_hbreak_req~q ),
	.prn(vcc));
defparam latched_oci_tb_hbreak_req.is_wysiwyg = "true";
defparam latched_oci_tb_hbreak_req.power_up = "low";

cyclonev_lcell_comb \F_iw~1 (
	.dataa(!hbreak_enabled1),
	.datab(!\latched_oci_tb_hbreak_req~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw~1 .extended_lut = "off";
defparam \F_iw~1 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \F_iw~1 .shared_arith = "off";

dffeas \D_iw[0] (
	.clk(clk_clk),
	.d(\F_iw[0]~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\F_iw~1_combout ),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\D_iw[0]~q ),
	.prn(vcc));
defparam \D_iw[0] .is_wysiwyg = "true";
defparam \D_iw[0] .power_up = "low";

cyclonev_lcell_comb \Equal4~2 (
	.dataa(!\D_iw[0]~q ),
	.datab(!\D_iw[1]~q ),
	.datac(!\D_iw[2]~q ),
	.datad(!\D_iw[3]~q ),
	.datae(!\D_iw[4]~q ),
	.dataf(!\D_iw[5]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal4~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal4~2 .extended_lut = "off";
defparam \Equal4~2 .lut_mask = 64'hFFEFFFFFFFFFFFFF;
defparam \Equal4~2 .shared_arith = "off";

cyclonev_lcell_comb \Equal4~3 (
	.dataa(!\D_iw[0]~q ),
	.datab(!\D_iw[1]~q ),
	.datac(!\D_iw[2]~q ),
	.datad(!\D_iw[3]~q ),
	.datae(!\D_iw[4]~q ),
	.dataf(!\D_iw[5]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal4~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal4~3 .extended_lut = "off";
defparam \Equal4~3 .lut_mask = 64'hEFFFFFFFFFFFFFFF;
defparam \Equal4~3 .shared_arith = "off";

cyclonev_lcell_comb \Equal4~4 (
	.dataa(!\D_iw[0]~q ),
	.datab(!\D_iw[1]~q ),
	.datac(!\D_iw[2]~q ),
	.datad(!\D_iw[3]~q ),
	.datae(!\D_iw[4]~q ),
	.dataf(!\D_iw[5]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal4~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal4~4 .extended_lut = "off";
defparam \Equal4~4 .lut_mask = 64'hFFFFEFFFFFFFFFFF;
defparam \Equal4~4 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_logic~0 (
	.dataa(!\D_iw[16]~q ),
	.datab(!\D_iw[11]~q ),
	.datac(!\D_ctrl_crst~0_combout ),
	.datad(!\Equal4~4_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_logic~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_logic~0 .extended_lut = "off";
defparam \D_ctrl_logic~0 .lut_mask = 64'hFFF7FFF7FFF7FFF7;
defparam \D_ctrl_logic~0 .shared_arith = "off";

cyclonev_lcell_comb D_ctrl_logic(
	.dataa(!\Equal4~2_combout ),
	.datab(!\Equal4~3_combout ),
	.datac(!\D_ctrl_logic~1_combout ),
	.datad(!\D_ctrl_logic~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_logic~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam D_ctrl_logic.extended_lut = "off";
defparam D_ctrl_logic.lut_mask = 64'hFF7FFF7FFF7FFF7F;
defparam D_ctrl_logic.shared_arith = "off";

dffeas E_ctrl_logic(
	.clk(clk_clk),
	.d(\D_ctrl_logic~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_ctrl_logic~q ),
	.prn(vcc));
defparam E_ctrl_logic.is_wysiwyg = "true";
defparam E_ctrl_logic.power_up = "low";

cyclonev_lcell_comb \E_wrctl_data_ienable_reg_irq16~0 (
	.dataa(!\E_ctrl_src2_choose_imm~q ),
	.datab(!\E_compare_op[1]~q ),
	.datac(!\E_compare_op[0]~q ),
	.datad(!\E_stw_data[16]~2_combout ),
	.datae(!\E_src2_imm[16]~q ),
	.dataf(!\E_src1[16]~9_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_wrctl_data_ienable_reg_irq16~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_wrctl_data_ienable_reg_irq16~0 .extended_lut = "off";
defparam \E_wrctl_data_ienable_reg_irq16~0 .lut_mask = 64'h6996966996696996;
defparam \E_wrctl_data_ienable_reg_irq16~0 .shared_arith = "off";

cyclonev_lcell_comb \D_control_reg_rddata_muxed[16]~0 (
	.dataa(!\D_iw[8]~q ),
	.datab(!\M_ipending_reg_irq16~q ),
	.datac(!\M_ienable_reg_irq16~q ),
	.datad(!\D_iw[7]~q ),
	.datae(!\D_iw[6]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_control_reg_rddata_muxed[16]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_control_reg_rddata_muxed[16]~0 .extended_lut = "off";
defparam \D_control_reg_rddata_muxed[16]~0 .lut_mask = 64'hBF7F7FBFBF7F7FBF;
defparam \D_control_reg_rddata_muxed[16]~0 .shared_arith = "off";

dffeas \E_control_reg_rddata[16] (
	.clk(clk_clk),
	.d(\D_control_reg_rddata_muxed[16]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_control_reg_rddata[16]~q ),
	.prn(vcc));
defparam \E_control_reg_rddata[16] .is_wysiwyg = "true";
defparam \E_control_reg_rddata[16] .power_up = "low";

cyclonev_lcell_comb \E_wrctl_data_ienable_reg_irq16~1 (
	.dataa(!\E_ctrl_retaddr~q ),
	.datab(!\E_ctrl_rdctl_inst~q ),
	.datac(!\E_control_reg_rddata[16]~q ),
	.datad(!\E_extra_pc[14]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_wrctl_data_ienable_reg_irq16~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_wrctl_data_ienable_reg_irq16~1 .extended_lut = "off";
defparam \E_wrctl_data_ienable_reg_irq16~1 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \E_wrctl_data_ienable_reg_irq16~1 .shared_arith = "off";

cyclonev_lcell_comb \E_wrctl_data_ienable_reg_irq16~2 (
	.dataa(!\E_ctrl_logic~q ),
	.datab(!\E_alu_result~0_combout ),
	.datac(!\Add8~13_sumout ),
	.datad(!\E_wrctl_data_ienable_reg_irq16~0_combout ),
	.datae(!\E_wrctl_data_ienable_reg_irq16~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_wrctl_data_ienable_reg_irq16~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_wrctl_data_ienable_reg_irq16~2 .extended_lut = "off";
defparam \E_wrctl_data_ienable_reg_irq16~2 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \E_wrctl_data_ienable_reg_irq16~2 .shared_arith = "off";

dffeas M_ienable_reg_irq16(
	.clk(clk_clk),
	.d(\E_wrctl_data_ienable_reg_irq16~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\M_ienable_reg_irq16~0_combout ),
	.q(\M_ienable_reg_irq16~q ),
	.prn(vcc));
defparam M_ienable_reg_irq16.is_wysiwyg = "true";
defparam M_ienable_reg_irq16.power_up = "low";

cyclonev_lcell_comb \M_ipending_reg_irq16_nxt~0 (
	.dataa(!\M_ienable_reg_irq16~q ),
	.datab(!\the_processor_cpu_nios2_oci|the_processor_cpu_nios2_avalon_reg|oci_ienable[16]~q ),
	.datac(!av_readdata_9),
	.datad(!av_readdata_8),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_ipending_reg_irq16_nxt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_ipending_reg_irq16_nxt~0 .extended_lut = "off";
defparam \M_ipending_reg_irq16_nxt~0 .lut_mask = 64'hDFFFDFFFDFFFDFFF;
defparam \M_ipending_reg_irq16_nxt~0 .shared_arith = "off";

dffeas M_ipending_reg_irq16(
	.clk(clk_clk),
	.d(\M_ipending_reg_irq16_nxt~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\M_ipending_reg_irq16~q ),
	.prn(vcc));
defparam M_ipending_reg_irq16.is_wysiwyg = "true";
defparam M_ipending_reg_irq16.power_up = "low";

cyclonev_lcell_comb \intr_req~0 (
	.dataa(!\M_ipending_reg_irq16~q ),
	.datab(!\M_status_reg_pie~q ),
	.datac(!\M_ipending_reg_irq1~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\intr_req~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \intr_req~0 .extended_lut = "off";
defparam \intr_req~0 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \intr_req~0 .shared_arith = "off";

cyclonev_lcell_comb \F_iw[24]~0 (
	.dataa(!\intr_req~0_combout ),
	.datab(!\processor_cpu_ic_data|the_altsyncram|auto_generated|q_b[24] ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[24]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[24]~0 .extended_lut = "off";
defparam \F_iw[24]~0 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \F_iw[24]~0 .shared_arith = "off";

dffeas \D_iw[24] (
	.clk(clk_clk),
	.d(\F_iw[24]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(\F_iw~1_combout ),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\D_iw[24]~q ),
	.prn(vcc));
defparam \D_iw[24] .is_wysiwyg = "true";
defparam \D_iw[24] .power_up = "low";

cyclonev_lcell_comb \D_dst_regnum[2]~1 (
	.dataa(!\D_iw[24]~q ),
	.datab(!\D_ctrl_b_not_src~0_combout ),
	.datac(!\D_iw[19]~q ),
	.datad(!\D_dst_regnum[4]~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_dst_regnum[2]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_dst_regnum[2]~1 .extended_lut = "off";
defparam \D_dst_regnum[2]~1 .lut_mask = 64'hDF1FDF1FDF1FDF1F;
defparam \D_dst_regnum[2]~1 .shared_arith = "off";

dffeas \E_dst_regnum[2] (
	.clk(clk_clk),
	.d(\D_dst_regnum[2]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_dst_regnum[2]~q ),
	.prn(vcc));
defparam \E_dst_regnum[2] .is_wysiwyg = "true";
defparam \E_dst_regnum[2] .power_up = "low";

cyclonev_lcell_comb \D_src2_hazard_E~0 (
	.dataa(!\E_dst_regnum[0]~q ),
	.datab(!\D_iw[22]~q ),
	.datac(!\E_dst_regnum[1]~q ),
	.datad(!\D_iw[23]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_hazard_E~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_hazard_E~0 .extended_lut = "off";
defparam \D_src2_hazard_E~0 .lut_mask = 64'h6996699669966996;
defparam \D_src2_hazard_E~0 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_hazard_E~1 (
	.dataa(!\E_dst_regnum[3]~q ),
	.datab(!\D_iw[25]~q ),
	.datac(!\E_dst_regnum[4]~q ),
	.datad(!\D_iw[26]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_hazard_E~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_hazard_E~1 .extended_lut = "off";
defparam \D_src2_hazard_E~1 .lut_mask = 64'h6996699669966996;
defparam \D_src2_hazard_E~1 .shared_arith = "off";

cyclonev_lcell_comb D_src2_hazard_E(
	.dataa(!\E_dst_regnum[2]~q ),
	.datab(!\D_iw[24]~q ),
	.datac(!\D_ctrl_b_not_src~0_combout ),
	.datad(!\E_wr_dst_reg~0_combout ),
	.datae(!\D_src2_hazard_E~0_combout ),
	.dataf(!\D_src2_hazard_E~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_hazard_E~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam D_src2_hazard_E.extended_lut = "off";
defparam D_src2_hazard_E.lut_mask = 64'hFF6FFFFFFFFFFFFF;
defparam D_src2_hazard_E.shared_arith = "off";

dffeas E_src2_hazard_M(
	.clk(clk_clk),
	.d(\D_src2_hazard_E~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_src2_hazard_M~q ),
	.prn(vcc));
defparam E_src2_hazard_M.is_wysiwyg = "true";
defparam E_src2_hazard_M.power_up = "low";

cyclonev_lcell_comb \E_stb_data[0]~0 (
	.dataa(!\E_src2_hazard_M~q ),
	.datab(!\M_shift_rot_result[0]~q ),
	.datac(!\M_ctrl_shift_rot~q ),
	.datad(!\av_ld_data_aligned_or_div[0]~q ),
	.datae(!\av_ld_or_div_done~q ),
	.dataf(!\M_alu_result[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_stb_data[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_stb_data[0]~0 .extended_lut = "off";
defparam \E_stb_data[0]~0 .lut_mask = 64'h7FFFF7FFFFFFFFFF;
defparam \E_stb_data[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \E_stb_data[0]~2 (
	.dataa(!\E_stb_data[0]~0_combout ),
	.datab(!\E_stb_data[0]~1_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_stb_data[0]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_stb_data[0]~2 .extended_lut = "off";
defparam \E_stb_data[0]~2 .lut_mask = 64'h7777777777777777;
defparam \E_stb_data[0]~2 .shared_arith = "off";

cyclonev_lcell_comb \Equal0~0 (
	.dataa(!\E_iw[4]~q ),
	.datab(!\E_iw[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~0 .extended_lut = "off";
defparam \Equal0~0 .lut_mask = 64'h7777777777777777;
defparam \Equal0~0 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_st~0 (
	.dataa(!\D_iw[0]~q ),
	.datab(!\D_iw[1]~q ),
	.datac(!\D_iw[2]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_st~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_st~0 .extended_lut = "off";
defparam \D_ctrl_st~0 .lut_mask = 64'hDFDFDFDFDFDFDFDF;
defparam \D_ctrl_st~0 .shared_arith = "off";

dffeas E_ctrl_st(
	.clk(clk_clk),
	.d(\D_ctrl_st~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\E_ctrl_st~q ),
	.prn(vcc));
defparam E_ctrl_st.is_wysiwyg = "true";
defparam E_ctrl_st.power_up = "low";

cyclonev_lcell_comb d_write_nxt(
	.dataa(!d_write1),
	.datab(!d_read1),
	.datac(!WideOr1),
	.datad(!read_accepted),
	.datae(!\E_ctrl_st~q ),
	.dataf(!\M_status_reg_pie~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d_write_nxt~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam d_write_nxt.extended_lut = "off";
defparam d_write_nxt.lut_mask = 64'hDF1FFFFFFFFFFFFF;
defparam d_write_nxt.shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[5]~1 (
	.dataa(!\E_ctrl_logic~q ),
	.datab(!\E_compare_op[1]~q ),
	.datac(!\E_compare_op[0]~q ),
	.datad(!\E_src1[5]~0_combout ),
	.datae(!\E_arith_src2[5]~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[5]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[5]~1 .extended_lut = "off";
defparam \E_alu_result[5]~1 .lut_mask = 64'h7DD7D77D7DD7D77D;
defparam \E_alu_result[5]~1 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[5]~2 (
	.dataa(!\E_ctrl_retaddr~q ),
	.datab(!\E_alu_result~0_combout ),
	.datac(!\E_extra_pc[3]~q ),
	.datad(!\Add8~1_sumout ),
	.datae(!\E_alu_result[5]~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[5]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[5]~2 .extended_lut = "off";
defparam \E_alu_result[5]~2 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \E_alu_result[5]~2 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[4]~3 (
	.dataa(!\E_ctrl_logic~q ),
	.datab(!\E_compare_op[1]~q ),
	.datac(!\E_compare_op[0]~q ),
	.datad(!\E_src1[4]~3_combout ),
	.datae(!\E_arith_src2[4]~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[4]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[4]~3 .extended_lut = "off";
defparam \E_alu_result[4]~3 .lut_mask = 64'h7DD7D77D7DD7D77D;
defparam \E_alu_result[4]~3 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[4]~4 (
	.dataa(!\E_ctrl_retaddr~q ),
	.datab(!\E_alu_result~0_combout ),
	.datac(!\E_extra_pc[2]~q ),
	.datad(!\Add8~5_sumout ),
	.datae(!\E_alu_result[4]~3_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[4]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[4]~4 .extended_lut = "off";
defparam \E_alu_result[4]~4 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \E_alu_result[4]~4 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[6]~64 (
	.dataa(!\E_src1[6]~6_combout ),
	.datab(!\E_compare_op[0]~q ),
	.datac(!\E_src2_imm[6]~q ),
	.datad(!\E_compare_op[1]~q ),
	.datae(!\E_ctrl_src2_choose_imm~q ),
	.dataf(!\E_ctrl_logic~q ),
	.datag(!\E_stb_data[6]~8_combout ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[6]~64_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[6]~64 .extended_lut = "on";
defparam \E_alu_result[6]~64 .lut_mask = 64'h6996699669966996;
defparam \E_alu_result[6]~64 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[6]~5 (
	.dataa(!\E_ctrl_retaddr~q ),
	.datab(!\E_alu_result~0_combout ),
	.datac(!\E_extra_pc[4]~q ),
	.datad(!\Add8~9_sumout ),
	.datae(!\E_alu_result[6]~64_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[6]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[6]~5 .extended_lut = "off";
defparam \E_alu_result[6]~5 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \E_alu_result[6]~5 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[15]~6 (
	.dataa(!\E_ctrl_logic~q ),
	.datab(!\E_compare_op[1]~q ),
	.datac(!\E_compare_op[0]~q ),
	.datad(!\E_src1[15]~10_combout ),
	.datae(!\E_arith_src2[15]~2_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[15]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[15]~6 .extended_lut = "off";
defparam \E_alu_result[15]~6 .lut_mask = 64'h7DD7D77D7DD7D77D;
defparam \E_alu_result[15]~6 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[15]~7 (
	.dataa(!\E_ctrl_retaddr~q ),
	.datab(!\E_alu_result~0_combout ),
	.datac(!\E_extra_pc[13]~q ),
	.datad(!\Add8~17_sumout ),
	.datae(!\E_alu_result[15]~6_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[15]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[15]~7 .extended_lut = "off";
defparam \E_alu_result[15]~7 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \E_alu_result[15]~7 .shared_arith = "off";

cyclonev_lcell_comb \E_arith_src2[14]~3 (
	.dataa(!\E_ctrl_src2_choose_imm~q ),
	.datab(!\E_stw_data[14]~4_combout ),
	.datac(!\E_src2_imm[14]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_arith_src2[14]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_arith_src2[14]~3 .extended_lut = "off";
defparam \E_arith_src2[14]~3 .lut_mask = 64'h2727272727272727;
defparam \E_arith_src2[14]~3 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[14]~8 (
	.dataa(!\E_ctrl_logic~q ),
	.datab(!\E_compare_op[1]~q ),
	.datac(!\E_compare_op[0]~q ),
	.datad(!\E_src1[14]~11_combout ),
	.datae(!\E_arith_src2[14]~3_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[14]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[14]~8 .extended_lut = "off";
defparam \E_alu_result[14]~8 .lut_mask = 64'h7DD7D77D7DD7D77D;
defparam \E_alu_result[14]~8 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[14]~9 (
	.dataa(!\E_ctrl_retaddr~q ),
	.datab(!\E_alu_result~0_combout ),
	.datac(!\E_extra_pc[12]~q ),
	.datad(!\Add8~21_sumout ),
	.datae(!\E_alu_result[14]~8_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[14]~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[14]~9 .extended_lut = "off";
defparam \E_alu_result[14]~9 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \E_alu_result[14]~9 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[13]~10 (
	.dataa(!\E_ctrl_logic~q ),
	.datab(!\E_compare_op[1]~q ),
	.datac(!\E_compare_op[0]~q ),
	.datad(!\E_src1[13]~12_combout ),
	.datae(!\E_arith_src2[13]~4_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[13]~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[13]~10 .extended_lut = "off";
defparam \E_alu_result[13]~10 .lut_mask = 64'h7DD7D77D7DD7D77D;
defparam \E_alu_result[13]~10 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[13]~11 (
	.dataa(!\E_ctrl_retaddr~q ),
	.datab(!\E_alu_result~0_combout ),
	.datac(!\E_extra_pc[11]~q ),
	.datad(!\Add8~25_sumout ),
	.datae(!\E_alu_result[13]~10_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[13]~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[13]~11 .extended_lut = "off";
defparam \E_alu_result[13]~11 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \E_alu_result[13]~11 .shared_arith = "off";

cyclonev_lcell_comb \E_arith_src2[12]~5 (
	.dataa(!\E_ctrl_src2_choose_imm~q ),
	.datab(!\E_stw_data[12]~5_combout ),
	.datac(!\E_src2_imm[12]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_arith_src2[12]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_arith_src2[12]~5 .extended_lut = "off";
defparam \E_arith_src2[12]~5 .lut_mask = 64'h2727272727272727;
defparam \E_arith_src2[12]~5 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[12]~12 (
	.dataa(!\E_ctrl_logic~q ),
	.datab(!\E_compare_op[1]~q ),
	.datac(!\E_compare_op[0]~q ),
	.datad(!\E_src1[12]~13_combout ),
	.datae(!\E_arith_src2[12]~5_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[12]~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[12]~12 .extended_lut = "off";
defparam \E_alu_result[12]~12 .lut_mask = 64'h7DD7D77D7DD7D77D;
defparam \E_alu_result[12]~12 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[12]~13 (
	.dataa(!\E_ctrl_retaddr~q ),
	.datab(!\E_alu_result~0_combout ),
	.datac(!\E_extra_pc[10]~q ),
	.datad(!\Add8~29_sumout ),
	.datae(!\E_alu_result[12]~12_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[12]~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[12]~13 .extended_lut = "off";
defparam \E_alu_result[12]~13 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \E_alu_result[12]~13 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[11]~14 (
	.dataa(!\E_ctrl_logic~q ),
	.datab(!\E_compare_op[1]~q ),
	.datac(!\E_compare_op[0]~q ),
	.datad(!\E_src1[11]~14_combout ),
	.datae(!\E_arith_src2[11]~6_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[11]~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[11]~14 .extended_lut = "off";
defparam \E_alu_result[11]~14 .lut_mask = 64'h7DD7D77D7DD7D77D;
defparam \E_alu_result[11]~14 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[11]~15 (
	.dataa(!\E_ctrl_retaddr~q ),
	.datab(!\E_alu_result~0_combout ),
	.datac(!\E_extra_pc[9]~q ),
	.datad(!\Add8~33_sumout ),
	.datae(!\E_alu_result[11]~14_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[11]~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[11]~15 .extended_lut = "off";
defparam \E_alu_result[11]~15 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \E_alu_result[11]~15 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[10]~60 (
	.dataa(!\E_src1[10]~17_combout ),
	.datab(!\E_compare_op[0]~q ),
	.datac(!\E_src2_imm[10]~q ),
	.datad(!\E_compare_op[1]~q ),
	.datae(!\E_ctrl_src2_choose_imm~q ),
	.dataf(!\E_ctrl_logic~q ),
	.datag(!\E_stw_data[10]~8_combout ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[10]~60_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[10]~60 .extended_lut = "on";
defparam \E_alu_result[10]~60 .lut_mask = 64'h6996699669966996;
defparam \E_alu_result[10]~60 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[10]~16 (
	.dataa(!\E_ctrl_retaddr~q ),
	.datab(!\E_alu_result~0_combout ),
	.datac(!\E_extra_pc[8]~q ),
	.datad(!\Add8~37_sumout ),
	.datae(!\E_alu_result[10]~60_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[10]~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[10]~16 .extended_lut = "off";
defparam \E_alu_result[10]~16 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \E_alu_result[10]~16 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[9]~17 (
	.dataa(!\E_ctrl_logic~q ),
	.datab(!\E_compare_op[1]~q ),
	.datac(!\E_compare_op[0]~q ),
	.datad(!\E_src1[9]~18_combout ),
	.datae(!\E_arith_src2[9]~7_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[9]~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[9]~17 .extended_lut = "off";
defparam \E_alu_result[9]~17 .lut_mask = 64'h7DD7D77D7DD7D77D;
defparam \E_alu_result[9]~17 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[9]~18 (
	.dataa(!\E_ctrl_retaddr~q ),
	.datab(!\E_alu_result~0_combout ),
	.datac(!\E_extra_pc[7]~q ),
	.datad(!\Add8~41_sumout ),
	.datae(!\E_alu_result[9]~17_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[9]~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[9]~18 .extended_lut = "off";
defparam \E_alu_result[9]~18 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \E_alu_result[9]~18 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[8]~56 (
	.dataa(!\E_src1[8]~21_combout ),
	.datab(!\E_compare_op[0]~q ),
	.datac(!\E_src2_imm[8]~q ),
	.datad(!\E_compare_op[1]~q ),
	.datae(!\E_ctrl_src2_choose_imm~q ),
	.dataf(!\E_ctrl_logic~q ),
	.datag(!\E_stw_data[8]~11_combout ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[8]~56_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[8]~56 .extended_lut = "on";
defparam \E_alu_result[8]~56 .lut_mask = 64'h6996699669966996;
defparam \E_alu_result[8]~56 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[8]~19 (
	.dataa(!\E_ctrl_retaddr~q ),
	.datab(!\E_alu_result~0_combout ),
	.datac(!\E_extra_pc[6]~q ),
	.datad(!\Add8~45_sumout ),
	.datae(!\E_alu_result[8]~56_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[8]~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[8]~19 .extended_lut = "off";
defparam \E_alu_result[8]~19 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \E_alu_result[8]~19 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[7]~20 (
	.dataa(!\E_ctrl_logic~q ),
	.datab(!\E_compare_op[1]~q ),
	.datac(!\E_compare_op[0]~q ),
	.datad(!\E_src1[7]~22_combout ),
	.datae(!\E_arith_src2[7]~8_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[7]~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[7]~20 .extended_lut = "off";
defparam \E_alu_result[7]~20 .lut_mask = 64'h7DD7D77D7DD7D77D;
defparam \E_alu_result[7]~20 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[7]~21 (
	.dataa(!\E_ctrl_retaddr~q ),
	.datab(!\E_alu_result~0_combout ),
	.datac(!\E_extra_pc[5]~q ),
	.datad(!\Add8~49_sumout ),
	.datae(!\E_alu_result[7]~20_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[7]~21_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[7]~21 .extended_lut = "off";
defparam \E_alu_result[7]~21 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \E_alu_result[7]~21 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[3]~22 (
	.dataa(!\E_ctrl_logic~q ),
	.datab(!\E_src1[3]~23_combout ),
	.datac(!\E_arith_src2[3]~9_combout ),
	.datad(!\E_compare_op[1]~q ),
	.datae(!\E_compare_op[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[3]~22_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[3]~22 .extended_lut = "off";
defparam \E_alu_result[3]~22 .lut_mask = 64'h7DD7D77D7DD7D77D;
defparam \E_alu_result[3]~22 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[3]~23 (
	.dataa(!\E_ctrl_retaddr~q ),
	.datab(!\E_extra_pc[1]~q ),
	.datac(!\Add8~53_sumout ),
	.datad(!\E_alu_result~0_combout ),
	.datae(!\E_alu_result[3]~22_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[3]~23_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[3]~23 .extended_lut = "off";
defparam \E_alu_result[3]~23 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \E_alu_result[3]~23 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[2]~24 (
	.dataa(!\E_ctrl_logic~q ),
	.datab(!\E_src1[2]~26_combout ),
	.datac(!\E_compare_op[1]~q ),
	.datad(!\E_compare_op[0]~q ),
	.datae(!\E_arith_src2[2]~10_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[2]~24_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[2]~24 .extended_lut = "off";
defparam \E_alu_result[2]~24 .lut_mask = 64'h7DD7D77D7DD7D77D;
defparam \E_alu_result[2]~24 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[2]~25 (
	.dataa(!\E_ctrl_retaddr~q ),
	.datab(!\E_alu_result~0_combout ),
	.datac(!\E_extra_pc[0]~q ),
	.datad(!\Add8~57_sumout ),
	.datae(!\E_alu_result[2]~24_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[2]~25_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[2]~25 .extended_lut = "off";
defparam \E_alu_result[2]~25 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \E_alu_result[2]~25 .shared_arith = "off";

cyclonev_lcell_comb d_read_nxt(
	.dataa(!d_read1),
	.datab(!WideOr1),
	.datac(!\M_status_reg_pie~0_combout ),
	.datad(!\E_ctrl_ld~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d_read_nxt~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam d_read_nxt.extended_lut = "off";
defparam d_read_nxt.lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam d_read_nxt.shared_arith = "off";

dffeas M_ctrl_break(
	.clk(clk_clk),
	.d(\E_ctrl_break~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\M_ctrl_break~q ),
	.prn(vcc));
defparam M_ctrl_break.is_wysiwyg = "true";
defparam M_ctrl_break.power_up = "low";

dffeas \M_iw[11] (
	.clk(clk_clk),
	.d(\E_iw[11]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\M_iw[11]~q ),
	.prn(vcc));
defparam \M_iw[11] .is_wysiwyg = "true";
defparam \M_iw[11] .power_up = "low";

dffeas \M_iw[1] (
	.clk(clk_clk),
	.d(\E_iw[1]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\M_iw[1]~q ),
	.prn(vcc));
defparam \M_iw[1] .is_wysiwyg = "true";
defparam \M_iw[1] .power_up = "low";

dffeas \M_iw[0] (
	.clk(clk_clk),
	.d(\E_iw[0]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\M_iw[0]~q ),
	.prn(vcc));
defparam \M_iw[0] .is_wysiwyg = "true";
defparam \M_iw[0] .power_up = "low";

dffeas \M_iw[16] (
	.clk(clk_clk),
	.d(\E_iw[16]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\M_iw[16]~q ),
	.prn(vcc));
defparam \M_iw[16] .is_wysiwyg = "true";
defparam \M_iw[16] .power_up = "low";

dffeas \M_iw[15] (
	.clk(clk_clk),
	.d(\E_iw[15]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\M_iw[15]~q ),
	.prn(vcc));
defparam \M_iw[15] .is_wysiwyg = "true";
defparam \M_iw[15] .power_up = "low";

dffeas \M_iw[14] (
	.clk(clk_clk),
	.d(\E_iw[14]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\M_iw[14]~q ),
	.prn(vcc));
defparam \M_iw[14] .is_wysiwyg = "true";
defparam \M_iw[14] .power_up = "low";

dffeas \M_iw[13] (
	.clk(clk_clk),
	.d(\E_iw[13]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\M_iw[13]~q ),
	.prn(vcc));
defparam \M_iw[13] .is_wysiwyg = "true";
defparam \M_iw[13] .power_up = "low";

dffeas \M_iw[12] (
	.clk(clk_clk),
	.d(\E_iw[12]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\M_iw[12]~q ),
	.prn(vcc));
defparam \M_iw[12] .is_wysiwyg = "true";
defparam \M_iw[12] .power_up = "low";

cyclonev_lcell_comb \hbreak_enabled~0 (
	.dataa(!\M_iw[16]~q ),
	.datab(!\M_iw[15]~q ),
	.datac(!\M_iw[14]~q ),
	.datad(!\M_iw[13]~q ),
	.datae(!\M_iw[12]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\hbreak_enabled~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \hbreak_enabled~0 .extended_lut = "off";
defparam \hbreak_enabled~0 .lut_mask = 64'hFFFFFFEFFFFFFFEF;
defparam \hbreak_enabled~0 .shared_arith = "off";

dffeas \M_iw[5] (
	.clk(clk_clk),
	.d(\E_iw[5]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\M_iw[5]~q ),
	.prn(vcc));
defparam \M_iw[5] .is_wysiwyg = "true";
defparam \M_iw[5] .power_up = "low";

dffeas \M_iw[2] (
	.clk(clk_clk),
	.d(\E_iw[2]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\M_iw[2]~q ),
	.prn(vcc));
defparam \M_iw[2] .is_wysiwyg = "true";
defparam \M_iw[2] .power_up = "low";

cyclonev_lcell_comb \hbreak_enabled~1 (
	.dataa(!\M_iw[4]~q ),
	.datab(!\M_iw[3]~q ),
	.datac(!\M_iw[5]~q ),
	.datad(!\M_iw[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\hbreak_enabled~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \hbreak_enabled~1 .extended_lut = "off";
defparam \hbreak_enabled~1 .lut_mask = 64'hFF7FFF7FFF7FFF7F;
defparam \hbreak_enabled~1 .shared_arith = "off";

cyclonev_lcell_comb \hbreak_enabled~2 (
	.dataa(!\M_iw[11]~q ),
	.datab(!\M_iw[1]~q ),
	.datac(!\M_iw[0]~q ),
	.datad(!\hbreak_enabled~0_combout ),
	.datae(!\hbreak_enabled~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\hbreak_enabled~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \hbreak_enabled~2 .extended_lut = "off";
defparam \hbreak_enabled~2 .lut_mask = 64'hF7FFFFFFF7FFFFFF;
defparam \hbreak_enabled~2 .shared_arith = "off";

cyclonev_lcell_comb \hbreak_enabled~3 (
	.dataa(!hbreak_enabled1),
	.datab(!\W_valid~0_combout ),
	.datac(!\M_ctrl_break~q ),
	.datad(!\hbreak_enabled~2_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\hbreak_enabled~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \hbreak_enabled~3 .extended_lut = "off";
defparam \hbreak_enabled~3 .lut_mask = 64'hDF1FDF1FDF1FDF1F;
defparam \hbreak_enabled~3 .shared_arith = "off";

cyclonev_lcell_comb \F_ic_fill_same_tag_line~0 (
	.dataa(!\F_pc[7]~q ),
	.datab(!\F_pc[6]~q ),
	.datac(!ic_fill_line_3),
	.datad(!ic_fill_line_4),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ic_fill_same_tag_line~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ic_fill_same_tag_line~0 .extended_lut = "off";
defparam \F_ic_fill_same_tag_line~0 .lut_mask = 64'h6996699669966996;
defparam \F_ic_fill_same_tag_line~0 .shared_arith = "off";

cyclonev_lcell_comb \F_ic_fill_same_tag_line~1 (
	.dataa(!\F_pc[3]~q ),
	.datab(!\F_pc[4]~q ),
	.datac(!ic_fill_line_0),
	.datad(!ic_fill_line_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ic_fill_same_tag_line~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ic_fill_same_tag_line~1 .extended_lut = "off";
defparam \F_ic_fill_same_tag_line~1 .lut_mask = 64'h6996699669966996;
defparam \F_ic_fill_same_tag_line~1 .shared_arith = "off";

cyclonev_lcell_comb \F_ic_fill_same_tag_line~2 (
	.dataa(!ic_fill_tag_1),
	.datab(!ic_fill_tag_0),
	.datac(!\F_pc[9]~q ),
	.datad(!\F_pc[10]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ic_fill_same_tag_line~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ic_fill_same_tag_line~2 .extended_lut = "off";
defparam \F_ic_fill_same_tag_line~2 .lut_mask = 64'h6996699669966996;
defparam \F_ic_fill_same_tag_line~2 .shared_arith = "off";

cyclonev_lcell_comb \F_ic_fill_same_tag_line~3 (
	.dataa(!ic_fill_tag_4),
	.datab(!ic_fill_tag_3),
	.datac(!\F_pc[12]~q ),
	.datad(!\F_pc[13]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ic_fill_same_tag_line~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ic_fill_same_tag_line~3 .extended_lut = "off";
defparam \F_ic_fill_same_tag_line~3 .lut_mask = 64'h6996699669966996;
defparam \F_ic_fill_same_tag_line~3 .shared_arith = "off";

cyclonev_lcell_comb \F_ic_fill_same_tag_line~4 (
	.dataa(!ic_fill_tag_5),
	.datab(!ic_fill_tag_2),
	.datac(!\F_pc[11]~q ),
	.datad(!\F_pc[14]~q ),
	.datae(!\F_ic_fill_same_tag_line~2_combout ),
	.dataf(!\F_ic_fill_same_tag_line~3_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ic_fill_same_tag_line~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ic_fill_same_tag_line~4 .extended_lut = "off";
defparam \F_ic_fill_same_tag_line~4 .lut_mask = 64'h6996FFFFFFFFFFFF;
defparam \F_ic_fill_same_tag_line~4 .shared_arith = "off";

cyclonev_lcell_comb \F_ic_fill_same_tag_line~5 (
	.dataa(!\F_pc[5]~q ),
	.datab(!ic_fill_line_2),
	.datac(!\F_ic_fill_same_tag_line~1_combout ),
	.datad(!\F_ic_fill_same_tag_line~4_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ic_fill_same_tag_line~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ic_fill_same_tag_line~5 .extended_lut = "off";
defparam \F_ic_fill_same_tag_line~5 .lut_mask = 64'h6FFF6FFF6FFF6FFF;
defparam \F_ic_fill_same_tag_line~5 .shared_arith = "off";

cyclonev_lcell_comb F_ic_fill_same_tag_line(
	.dataa(!ic_fill_line_5),
	.datab(!\F_pc[8]~q ),
	.datac(!\F_ic_fill_same_tag_line~0_combout ),
	.datad(!\F_ic_fill_same_tag_line~5_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ic_fill_same_tag_line~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam F_ic_fill_same_tag_line.extended_lut = "off";
defparam F_ic_fill_same_tag_line.lut_mask = 64'h6FFF6FFF6FFF6FFF;
defparam F_ic_fill_same_tag_line.shared_arith = "off";

dffeas D_ic_fill_same_tag_line(
	.clk(clk_clk),
	.d(\F_ic_fill_same_tag_line~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\D_ic_fill_same_tag_line~q ),
	.prn(vcc));
defparam D_ic_fill_same_tag_line.is_wysiwyg = "true";
defparam D_ic_fill_same_tag_line.power_up = "low";

cyclonev_lcell_comb \E_ctrl_invalidate_i~0 (
	.dataa(!\E_iw[16]~q ),
	.datab(!\E_iw[15]~q ),
	.datac(!\E_iw[13]~q ),
	.datad(!\E_iw[12]~q ),
	.datae(!\E_iw[11]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_ctrl_invalidate_i~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_ctrl_invalidate_i~0 .extended_lut = "off";
defparam \E_ctrl_invalidate_i~0 .lut_mask = 64'h9669699696696996;
defparam \E_ctrl_invalidate_i~0 .shared_arith = "off";

cyclonev_lcell_comb \E_ctrl_invalidate_i~1 (
	.dataa(!\E_iw[14]~q ),
	.datab(!\Equal130~0_combout ),
	.datac(!\E_ctrl_invalidate_i~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_ctrl_invalidate_i~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_ctrl_invalidate_i~1 .extended_lut = "off";
defparam \E_ctrl_invalidate_i~1 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \E_ctrl_invalidate_i~1 .shared_arith = "off";

dffeas M_ctrl_invalidate_i(
	.clk(clk_clk),
	.d(\E_ctrl_invalidate_i~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\W_stall~combout ),
	.q(\M_ctrl_invalidate_i~q ),
	.prn(vcc));
defparam M_ctrl_invalidate_i.is_wysiwyg = "true";
defparam M_ctrl_invalidate_i.power_up = "low";

cyclonev_lcell_comb ic_fill_prevent_refill_nxt(
	.dataa(!\M_valid_from_E~q ),
	.datab(!\ic_fill_prevent_refill~q ),
	.datac(!\D_ic_fill_starting~0_combout ),
	.datad(!\M_ctrl_invalidate_i~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_fill_prevent_refill_nxt~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam ic_fill_prevent_refill_nxt.extended_lut = "off";
defparam ic_fill_prevent_refill_nxt.lut_mask = 64'hFFBFFFBFFFBFFFBF;
defparam ic_fill_prevent_refill_nxt.shared_arith = "off";

dffeas ic_fill_prevent_refill(
	.clk(clk_clk),
	.d(\ic_fill_prevent_refill_nxt~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ic_fill_prevent_refill~q ),
	.prn(vcc));
defparam ic_fill_prevent_refill.is_wysiwyg = "true";
defparam ic_fill_prevent_refill.power_up = "low";

cyclonev_lcell_comb \D_ic_fill_starting~0 (
	.dataa(!\M_pipe_flush~q ),
	.datab(!\D_ic_fill_same_tag_line~q ),
	.datac(!\ic_fill_prevent_refill~q ),
	.datad(!\ic_fill_active~q ),
	.datae(!\D_iw_valid~q ),
	.dataf(!\D_kill~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ic_fill_starting~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ic_fill_starting~0 .extended_lut = "off";
defparam \D_ic_fill_starting~0 .lut_mask = 64'hFFFFFFFFFFFFFFFD;
defparam \D_ic_fill_starting~0 .shared_arith = "off";

dffeas \ic_fill_initial_offset[2] (
	.clk(clk_clk),
	.d(\D_pc[2]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\D_ic_fill_starting~0_combout ),
	.q(\ic_fill_initial_offset[2]~q ),
	.prn(vcc));
defparam \ic_fill_initial_offset[2] .is_wysiwyg = "true";
defparam \ic_fill_initial_offset[2] .power_up = "low";

dffeas \ic_fill_initial_offset[0] (
	.clk(clk_clk),
	.d(\D_pc[0]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\D_ic_fill_starting~0_combout ),
	.q(\ic_fill_initial_offset[0]~q ),
	.prn(vcc));
defparam \ic_fill_initial_offset[0] .is_wysiwyg = "true";
defparam \ic_fill_initial_offset[0] .power_up = "low";

dffeas D_ic_fill_starting_d1(
	.clk(clk_clk),
	.d(\D_ic_fill_starting~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\D_ic_fill_starting_d1~q ),
	.prn(vcc));
defparam D_ic_fill_starting_d1.is_wysiwyg = "true";
defparam D_ic_fill_starting_d1.power_up = "low";

cyclonev_lcell_comb \ic_fill_dp_offset_nxt[0]~1 (
	.dataa(!\ic_fill_dp_offset[0]~q ),
	.datab(!\ic_fill_initial_offset[0]~q ),
	.datac(!\D_ic_fill_starting_d1~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_fill_dp_offset_nxt[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_fill_dp_offset_nxt[0]~1 .extended_lut = "off";
defparam \ic_fill_dp_offset_nxt[0]~1 .lut_mask = 64'hA3A3A3A3A3A3A3A3;
defparam \ic_fill_dp_offset_nxt[0]~1 .shared_arith = "off";

dffeas i_readdatavalid_d1(
	.clk(clk_clk),
	.d(WideOr11),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_readdatavalid_d1~q ),
	.prn(vcc));
defparam i_readdatavalid_d1.is_wysiwyg = "true";
defparam i_readdatavalid_d1.power_up = "low";

cyclonev_lcell_comb \ic_fill_dp_offset_en~0 (
	.dataa(!\i_readdatavalid_d1~q ),
	.datab(!\D_ic_fill_starting_d1~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_fill_dp_offset_en~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_fill_dp_offset_en~0 .extended_lut = "off";
defparam \ic_fill_dp_offset_en~0 .lut_mask = 64'h7777777777777777;
defparam \ic_fill_dp_offset_en~0 .shared_arith = "off";

dffeas \ic_fill_dp_offset[0] (
	.clk(clk_clk),
	.d(\ic_fill_dp_offset_nxt[0]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ic_fill_dp_offset_en~0_combout ),
	.q(\ic_fill_dp_offset[0]~q ),
	.prn(vcc));
defparam \ic_fill_dp_offset[0] .is_wysiwyg = "true";
defparam \ic_fill_dp_offset[0] .power_up = "low";

dffeas \ic_fill_initial_offset[1] (
	.clk(clk_clk),
	.d(\D_pc[1]~q ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\D_ic_fill_starting~0_combout ),
	.q(\ic_fill_initial_offset[1]~q ),
	.prn(vcc));
defparam \ic_fill_initial_offset[1] .is_wysiwyg = "true";
defparam \ic_fill_initial_offset[1] .power_up = "low";

cyclonev_lcell_comb \ic_fill_dp_offset_nxt[1]~2 (
	.dataa(!\ic_fill_dp_offset[0]~q ),
	.datab(!\ic_fill_dp_offset[1]~q ),
	.datac(!\D_ic_fill_starting_d1~q ),
	.datad(!\ic_fill_initial_offset[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_fill_dp_offset_nxt[1]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_fill_dp_offset_nxt[1]~2 .extended_lut = "off";
defparam \ic_fill_dp_offset_nxt[1]~2 .lut_mask = 64'h96FF96FF96FF96FF;
defparam \ic_fill_dp_offset_nxt[1]~2 .shared_arith = "off";

dffeas \ic_fill_dp_offset[1] (
	.clk(clk_clk),
	.d(\ic_fill_dp_offset_nxt[1]~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ic_fill_dp_offset_en~0_combout ),
	.q(\ic_fill_dp_offset[1]~q ),
	.prn(vcc));
defparam \ic_fill_dp_offset[1] .is_wysiwyg = "true";
defparam \ic_fill_dp_offset[1] .power_up = "low";

dffeas \ic_fill_dp_offset[2] (
	.clk(clk_clk),
	.d(\ic_fill_dp_offset_nxt[2]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ic_fill_dp_offset_en~0_combout ),
	.q(\ic_fill_dp_offset[2]~q ),
	.prn(vcc));
defparam \ic_fill_dp_offset[2] .is_wysiwyg = "true";
defparam \ic_fill_dp_offset[2] .power_up = "low";

cyclonev_lcell_comb \ic_fill_dp_offset_nxt[2]~0 (
	.dataa(!\ic_fill_dp_offset[0]~q ),
	.datab(!\ic_fill_dp_offset[1]~q ),
	.datac(!\ic_fill_dp_offset[2]~q ),
	.datad(!\D_ic_fill_starting_d1~q ),
	.datae(!\ic_fill_initial_offset[2]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_fill_dp_offset_nxt[2]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_fill_dp_offset_nxt[2]~0 .extended_lut = "off";
defparam \ic_fill_dp_offset_nxt[2]~0 .lut_mask = 64'h6996FFFF6996FFFF;
defparam \ic_fill_dp_offset_nxt[2]~0 .shared_arith = "off";

cyclonev_lcell_comb \ic_fill_active_nxt~0 (
	.dataa(!\i_readdatavalid_d1~q ),
	.datab(!\ic_fill_initial_offset[0]~q ),
	.datac(!\ic_fill_dp_offset_nxt[0]~1_combout ),
	.datad(!\ic_fill_initial_offset[1]~q ),
	.datae(!\ic_fill_dp_offset_nxt[1]~2_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_fill_active_nxt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_fill_active_nxt~0 .extended_lut = "off";
defparam \ic_fill_active_nxt~0 .lut_mask = 64'h7DD7D77D7DD7D77D;
defparam \ic_fill_active_nxt~0 .shared_arith = "off";

cyclonev_lcell_comb \ic_fill_active_nxt~1 (
	.dataa(!\ic_fill_active~q ),
	.datab(!\D_ic_fill_starting~0_combout ),
	.datac(!\ic_fill_initial_offset[2]~q ),
	.datad(!\ic_fill_dp_offset_nxt[2]~0_combout ),
	.datae(!\ic_fill_active_nxt~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_fill_active_nxt~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_fill_active_nxt~1 .extended_lut = "off";
defparam \ic_fill_active_nxt~1 .lut_mask = 64'hFFFF7FF7FFFF7FF7;
defparam \ic_fill_active_nxt~1 .shared_arith = "off";

dffeas ic_fill_active(
	.clk(clk_clk),
	.d(\ic_fill_active_nxt~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ic_fill_active~q ),
	.prn(vcc));
defparam ic_fill_active.is_wysiwyg = "true";
defparam ic_fill_active.power_up = "low";

cyclonev_lcell_comb \ic_fill_ap_cnt_nxt[0]~3 (
	.dataa(!nonposted_cmd_accepted),
	.datab(!\ic_fill_ap_cnt[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_fill_ap_cnt_nxt[0]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_fill_ap_cnt_nxt[0]~3 .extended_lut = "off";
defparam \ic_fill_ap_cnt_nxt[0]~3 .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \ic_fill_ap_cnt_nxt[0]~3 .shared_arith = "off";

cyclonev_lcell_comb \ic_fill_ap_cnt[2]~0 (
	.dataa(!nonposted_cmd_accepted),
	.datab(!\D_ic_fill_starting~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_fill_ap_cnt[2]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_fill_ap_cnt[2]~0 .extended_lut = "off";
defparam \ic_fill_ap_cnt[2]~0 .lut_mask = 64'h7777777777777777;
defparam \ic_fill_ap_cnt[2]~0 .shared_arith = "off";

dffeas \ic_fill_ap_cnt[0] (
	.clk(clk_clk),
	.d(\ic_fill_ap_cnt_nxt[0]~3_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ic_fill_ap_cnt[2]~0_combout ),
	.q(\ic_fill_ap_cnt[0]~q ),
	.prn(vcc));
defparam \ic_fill_ap_cnt[0] .is_wysiwyg = "true";
defparam \ic_fill_ap_cnt[0] .power_up = "low";

cyclonev_lcell_comb \ic_fill_ap_cnt_nxt[1]~2 (
	.dataa(!nonposted_cmd_accepted),
	.datab(!\ic_fill_ap_cnt[1]~q ),
	.datac(!\ic_fill_ap_cnt[0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_fill_ap_cnt_nxt[1]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_fill_ap_cnt_nxt[1]~2 .extended_lut = "off";
defparam \ic_fill_ap_cnt_nxt[1]~2 .lut_mask = 64'h7D7D7D7D7D7D7D7D;
defparam \ic_fill_ap_cnt_nxt[1]~2 .shared_arith = "off";

dffeas \ic_fill_ap_cnt[1] (
	.clk(clk_clk),
	.d(\ic_fill_ap_cnt_nxt[1]~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ic_fill_ap_cnt[2]~0_combout ),
	.q(\ic_fill_ap_cnt[1]~q ),
	.prn(vcc));
defparam \ic_fill_ap_cnt[1] .is_wysiwyg = "true";
defparam \ic_fill_ap_cnt[1] .power_up = "low";

cyclonev_lcell_comb \ic_fill_ap_cnt_nxt[2]~1 (
	.dataa(!nonposted_cmd_accepted),
	.datab(!\ic_fill_ap_cnt[2]~q ),
	.datac(!\ic_fill_ap_cnt[1]~q ),
	.datad(!\ic_fill_ap_cnt[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_fill_ap_cnt_nxt[2]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_fill_ap_cnt_nxt[2]~1 .extended_lut = "off";
defparam \ic_fill_ap_cnt_nxt[2]~1 .lut_mask = 64'hD77DD77DD77DD77D;
defparam \ic_fill_ap_cnt_nxt[2]~1 .shared_arith = "off";

dffeas \ic_fill_ap_cnt[2] (
	.clk(clk_clk),
	.d(\ic_fill_ap_cnt_nxt[2]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ic_fill_ap_cnt[2]~0_combout ),
	.q(\ic_fill_ap_cnt[2]~q ),
	.prn(vcc));
defparam \ic_fill_ap_cnt[2] .is_wysiwyg = "true";
defparam \ic_fill_ap_cnt[2] .power_up = "low";

cyclonev_lcell_comb \ic_fill_ap_cnt_nxt[3]~0 (
	.dataa(!nonposted_cmd_accepted),
	.datab(!\ic_fill_ap_cnt[3]~q ),
	.datac(!\ic_fill_ap_cnt[2]~q ),
	.datad(!\ic_fill_ap_cnt[1]~q ),
	.datae(!\ic_fill_ap_cnt[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_fill_ap_cnt_nxt[3]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_fill_ap_cnt_nxt[3]~0 .extended_lut = "off";
defparam \ic_fill_ap_cnt_nxt[3]~0 .lut_mask = 64'h7DD7D77D7DD7D77D;
defparam \ic_fill_ap_cnt_nxt[3]~0 .shared_arith = "off";

dffeas \ic_fill_ap_cnt[3] (
	.clk(clk_clk),
	.d(\ic_fill_ap_cnt_nxt[3]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ic_fill_ap_cnt[2]~0_combout ),
	.q(\ic_fill_ap_cnt[3]~q ),
	.prn(vcc));
defparam \ic_fill_ap_cnt[3] .is_wysiwyg = "true";
defparam \ic_fill_ap_cnt[3] .power_up = "low";

cyclonev_lcell_comb \i_read_nxt~0 (
	.dataa(!clr_break_line1),
	.datab(!WideOr0),
	.datac(!\ic_fill_active~q ),
	.datad(!\ic_fill_ap_cnt[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\i_read_nxt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \i_read_nxt~0 .extended_lut = "off";
defparam \i_read_nxt~0 .lut_mask = 64'hF7FFF7FFF7FFF7FF;
defparam \i_read_nxt~0 .shared_arith = "off";

cyclonev_lcell_comb \i_read_nxt~1 (
	.dataa(!has_pending_responses),
	.datab(!i_read1),
	.datac(!Equal1),
	.datad(!last_dest_id_1),
	.datae(!\i_read_nxt~0_combout ),
	.dataf(!\D_ic_fill_starting~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\i_read_nxt~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \i_read_nxt~1 .extended_lut = "off";
defparam \i_read_nxt~1 .lut_mask = 64'hFFFF7FF7FFFFFFFF;
defparam \i_read_nxt~1 .shared_arith = "off";

cyclonev_lcell_comb \ic_tag_wraddress_nxt~0 (
	.dataa(!\D_ic_fill_starting~0_combout ),
	.datab(!ic_fill_line_5),
	.datac(!\D_pc[8]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_tag_wraddress_nxt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_tag_wraddress_nxt~0 .extended_lut = "off";
defparam \ic_tag_wraddress_nxt~0 .lut_mask = 64'h2727272727272727;
defparam \ic_tag_wraddress_nxt~0 .shared_arith = "off";

cyclonev_lcell_comb \ic_tag_wraddress_nxt~1 (
	.dataa(!\D_ic_fill_starting~0_combout ),
	.datab(!ic_fill_line_0),
	.datac(!\D_pc[3]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_tag_wraddress_nxt~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_tag_wraddress_nxt~1 .extended_lut = "off";
defparam \ic_tag_wraddress_nxt~1 .lut_mask = 64'h2727272727272727;
defparam \ic_tag_wraddress_nxt~1 .shared_arith = "off";

cyclonev_lcell_comb \ic_tag_wraddress_nxt~2 (
	.dataa(!\D_ic_fill_starting~0_combout ),
	.datab(!ic_fill_line_1),
	.datac(!\D_pc[4]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_tag_wraddress_nxt~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_tag_wraddress_nxt~2 .extended_lut = "off";
defparam \ic_tag_wraddress_nxt~2 .lut_mask = 64'h2727272727272727;
defparam \ic_tag_wraddress_nxt~2 .shared_arith = "off";

cyclonev_lcell_comb \ic_tag_wraddress_nxt~3 (
	.dataa(!\D_ic_fill_starting~0_combout ),
	.datab(!ic_fill_line_2),
	.datac(!\D_pc[5]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_tag_wraddress_nxt~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_tag_wraddress_nxt~3 .extended_lut = "off";
defparam \ic_tag_wraddress_nxt~3 .lut_mask = 64'h2727272727272727;
defparam \ic_tag_wraddress_nxt~3 .shared_arith = "off";

cyclonev_lcell_comb \ic_tag_wraddress_nxt~4 (
	.dataa(!\D_ic_fill_starting~0_combout ),
	.datab(!ic_fill_line_3),
	.datac(!\D_pc[6]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_tag_wraddress_nxt~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_tag_wraddress_nxt~4 .extended_lut = "off";
defparam \ic_tag_wraddress_nxt~4 .lut_mask = 64'h2727272727272727;
defparam \ic_tag_wraddress_nxt~4 .shared_arith = "off";

cyclonev_lcell_comb \ic_tag_wraddress_nxt~5 (
	.dataa(!\D_ic_fill_starting~0_combout ),
	.datab(!ic_fill_line_4),
	.datac(!\D_pc[7]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_tag_wraddress_nxt~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_tag_wraddress_nxt~5 .extended_lut = "off";
defparam \ic_tag_wraddress_nxt~5 .lut_mask = 64'h2727272727272727;
defparam \ic_tag_wraddress_nxt~5 .shared_arith = "off";

cyclonev_lcell_comb \ic_fill_ap_offset_nxt[0]~0 (
	.dataa(!nonposted_cmd_accepted),
	.datab(!\D_pc[0]~q ),
	.datac(!ic_fill_ap_offset_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_fill_ap_offset_nxt[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_fill_ap_offset_nxt[0]~0 .extended_lut = "off";
defparam \ic_fill_ap_offset_nxt[0]~0 .lut_mask = 64'hB1B1B1B1B1B1B1B1;
defparam \ic_fill_ap_offset_nxt[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \ic_fill_ap_offset_nxt[1]~1 (
	.dataa(!nonposted_cmd_accepted),
	.datab(!\D_pc[1]~q ),
	.datac(!ic_fill_ap_offset_0),
	.datad(!ic_fill_ap_offset_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_fill_ap_offset_nxt[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_fill_ap_offset_nxt[1]~1 .extended_lut = "off";
defparam \ic_fill_ap_offset_nxt[1]~1 .lut_mask = 64'hB77BB77BB77BB77B;
defparam \ic_fill_ap_offset_nxt[1]~1 .shared_arith = "off";

cyclonev_lcell_comb \ic_fill_ap_offset_nxt[2]~2 (
	.dataa(!nonposted_cmd_accepted),
	.datab(!\D_pc[2]~q ),
	.datac(!ic_fill_ap_offset_0),
	.datad(!ic_fill_ap_offset_1),
	.datae(!ic_fill_ap_offset_2),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_fill_ap_offset_nxt[2]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_fill_ap_offset_nxt[2]~2 .extended_lut = "off";
defparam \ic_fill_ap_offset_nxt[2]~2 .lut_mask = 64'h7BB7B77B7BB7B77B;
defparam \ic_fill_ap_offset_nxt[2]~2 .shared_arith = "off";

cyclonev_lcell_comb \E_mem_byte_en~0 (
	.dataa(!\E_iw[4]~q ),
	.datab(!\E_iw[3]~q ),
	.datac(!\Add8~65_sumout ),
	.datad(!\Add8~69_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_mem_byte_en~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_mem_byte_en~0 .extended_lut = "off";
defparam \E_mem_byte_en~0 .lut_mask = 64'hFFF7FFF7FFF7FFF7;
defparam \E_mem_byte_en~0 .shared_arith = "off";

cyclonev_lcell_comb \E_mem_byte_en[2]~1 (
	.dataa(!\E_iw[4]~q ),
	.datab(!\E_iw[3]~q ),
	.datac(!\Add8~65_sumout ),
	.datad(!\Add8~69_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_mem_byte_en[2]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_mem_byte_en[2]~1 .extended_lut = "off";
defparam \E_mem_byte_en[2]~1 .lut_mask = 64'hF7FFF7FFF7FFF7FF;
defparam \E_mem_byte_en[2]~1 .shared_arith = "off";

cyclonev_lcell_comb \E_mem_byte_en[1]~2 (
	.dataa(!\E_iw[4]~q ),
	.datab(!\E_iw[3]~q ),
	.datac(!\Add8~65_sumout ),
	.datad(!\Add8~69_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_mem_byte_en[1]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_mem_byte_en[1]~2 .extended_lut = "off";
defparam \E_mem_byte_en[1]~2 .lut_mask = 64'hFF7FFF7FFF7FFF7F;
defparam \E_mem_byte_en[1]~2 .shared_arith = "off";

cyclonev_lcell_comb \E_st_data[24]~0 (
	.dataa(!\E_stb_data[0]~2_combout ),
	.datab(!\E_iw[4]~q ),
	.datac(!\E_iw[3]~q ),
	.datad(!\E_stw_data[8]~11_combout ),
	.datae(!\E_stw_data[24]~20_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_st_data[24]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_st_data[24]~0 .extended_lut = "off";
defparam \E_st_data[24]~0 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \E_st_data[24]~0 .shared_arith = "off";

cyclonev_lcell_comb \E_mem_byte_en[3]~3 (
	.dataa(!\E_iw[4]~q ),
	.datab(!\E_iw[3]~q ),
	.datac(!\Add8~65_sumout ),
	.datad(!\Add8~69_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_mem_byte_en[3]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_mem_byte_en[3]~3 .extended_lut = "off";
defparam \E_mem_byte_en[3]~3 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \E_mem_byte_en[3]~3 .shared_arith = "off";

cyclonev_lcell_comb \E_st_data[29]~1 (
	.dataa(!\E_iw[4]~q ),
	.datab(!\E_iw[3]~q ),
	.datac(!\E_stb_data[5]~14_combout ),
	.datad(!\E_stw_data[13]~13_combout ),
	.datae(!\E_stw_data[29]~22_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_st_data[29]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_st_data[29]~1 .extended_lut = "off";
defparam \E_st_data[29]~1 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \E_st_data[29]~1 .shared_arith = "off";

cyclonev_lcell_comb \E_st_data[28]~2 (
	.dataa(!\E_iw[4]~q ),
	.datab(!\E_iw[3]~q ),
	.datac(!\E_stb_data[4]~5_combout ),
	.datad(!\E_stw_data[12]~5_combout ),
	.datae(!\E_stw_data[28]~28_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_st_data[28]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_st_data[28]~2 .extended_lut = "off";
defparam \E_st_data[28]~2 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \E_st_data[28]~2 .shared_arith = "off";

cyclonev_lcell_comb \E_st_data[30]~3 (
	.dataa(!\E_iw[4]~q ),
	.datab(!\E_iw[3]~q ),
	.datac(!\E_stb_data[6]~8_combout ),
	.datad(!\E_stw_data[14]~4_combout ),
	.datae(!\E_stw_data[30]~17_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_st_data[30]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_st_data[30]~3 .extended_lut = "off";
defparam \E_st_data[30]~3 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \E_st_data[30]~3 .shared_arith = "off";

cyclonev_lcell_comb \E_st_data[31]~4 (
	.dataa(!\E_src2_hazard_M~q ),
	.datab(!\M_wr_data_unfiltered[31]~17_combout ),
	.datac(!\E_src2_prelim[31]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_st_data[31]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_st_data[31]~4 .extended_lut = "off";
defparam \E_st_data[31]~4 .lut_mask = 64'h2727272727272727;
defparam \E_st_data[31]~4 .shared_arith = "off";

cyclonev_lcell_comb \E_st_data[31]~5 (
	.dataa(!\E_iw[4]~q ),
	.datab(!\E_iw[3]~q ),
	.datac(!\E_stb_data[7]~15_combout ),
	.datad(!\E_stw_data[15]~3_combout ),
	.datae(!\E_st_data[31]~4_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_st_data[31]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_st_data[31]~5 .extended_lut = "off";
defparam \E_st_data[31]~5 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \E_st_data[31]~5 .shared_arith = "off";

cyclonev_lcell_comb \E_st_data[27]~6 (
	.dataa(!\E_stb_data[3]~13_combout ),
	.datab(!\E_iw[4]~q ),
	.datac(!\E_iw[3]~q ),
	.datad(!\E_stw_data[11]~14_combout ),
	.datae(!\E_stw_data[27]~37_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_st_data[27]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_st_data[27]~6 .extended_lut = "off";
defparam \E_st_data[27]~6 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \E_st_data[27]~6 .shared_arith = "off";

cyclonev_lcell_comb \E_st_data[26]~7 (
	.dataa(!\E_stb_data[2]~11_combout ),
	.datab(!\E_iw[4]~q ),
	.datac(!\E_iw[3]~q ),
	.datad(!\E_stw_data[10]~8_combout ),
	.datae(!\E_stw_data[26]~40_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_st_data[26]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_st_data[26]~7 .extended_lut = "off";
defparam \E_st_data[26]~7 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \E_st_data[26]~7 .shared_arith = "off";

cyclonev_lcell_comb \E_st_data[25]~8 (
	.dataa(!\E_stb_data[1]~12_combout ),
	.datab(!\E_iw[4]~q ),
	.datac(!\E_iw[3]~q ),
	.datad(!\E_stw_data[9]~12_combout ),
	.datae(!\E_stw_data[25]~41_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_st_data[25]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_st_data[25]~8 .extended_lut = "off";
defparam \E_st_data[25]~8 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \E_st_data[25]~8 .shared_arith = "off";

endmodule

module processor_processor_cpu_ic_data_module (
	q_b_24,
	q_b_0,
	q_b_1,
	q_b_2,
	q_b_3,
	q_b_4,
	q_b_5,
	q_b_22,
	q_b_23,
	q_b_25,
	q_b_26,
	q_b_14,
	q_b_12,
	q_b_11,
	q_b_16,
	q_b_15,
	q_b_13,
	q_b_21,
	q_b_29,
	q_b_27,
	q_b_28,
	q_b_30,
	q_b_31,
	q_b_10,
	q_b_6,
	q_b_8,
	q_b_7,
	q_b_20,
	q_b_19,
	q_b_18,
	q_b_17,
	q_b_9,
	W_stall,
	ic_fill_line_5,
	i_readdatavalid_d1,
	i_readdata_d1_24,
	ic_fill_dp_offset_0,
	ic_fill_dp_offset_1,
	ic_fill_dp_offset_2,
	ic_fill_line_0,
	ic_fill_line_1,
	ic_fill_line_2,
	ic_fill_line_3,
	ic_fill_line_4,
	F_ic_data_rd_addr_nxt_0,
	F_ic_data_rd_addr_nxt_1,
	F_ic_data_rd_addr_nxt_2,
	F_ic_tag_rd_addr_nxt_0,
	F_ic_tag_rd_addr_nxt_1,
	F_ic_tag_rd_addr_nxt_2,
	F_ic_tag_rd_addr_nxt_3,
	F_ic_tag_rd_addr_nxt_4,
	F_ic_tag_rd_addr_nxt_5,
	i_readdata_d1_0,
	i_readdata_d1_1,
	i_readdata_d1_2,
	i_readdata_d1_3,
	i_readdata_d1_4,
	i_readdata_d1_5,
	i_readdata_d1_22,
	i_readdata_d1_23,
	i_readdata_d1_25,
	i_readdata_d1_26,
	i_readdata_d1_14,
	i_readdata_d1_12,
	i_readdata_d1_11,
	i_readdata_d1_16,
	i_readdata_d1_15,
	i_readdata_d1_13,
	i_readdata_d1_21,
	i_readdata_d1_29,
	i_readdata_d1_27,
	i_readdata_d1_28,
	i_readdata_d1_30,
	i_readdata_d1_31,
	i_readdata_d1_10,
	i_readdata_d1_6,
	i_readdata_d1_8,
	i_readdata_d1_7,
	i_readdata_d1_20,
	i_readdata_d1_19,
	i_readdata_d1_18,
	i_readdata_d1_17,
	i_readdata_d1_9,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_24;
output 	q_b_0;
output 	q_b_1;
output 	q_b_2;
output 	q_b_3;
output 	q_b_4;
output 	q_b_5;
output 	q_b_22;
output 	q_b_23;
output 	q_b_25;
output 	q_b_26;
output 	q_b_14;
output 	q_b_12;
output 	q_b_11;
output 	q_b_16;
output 	q_b_15;
output 	q_b_13;
output 	q_b_21;
output 	q_b_29;
output 	q_b_27;
output 	q_b_28;
output 	q_b_30;
output 	q_b_31;
output 	q_b_10;
output 	q_b_6;
output 	q_b_8;
output 	q_b_7;
output 	q_b_20;
output 	q_b_19;
output 	q_b_18;
output 	q_b_17;
output 	q_b_9;
input 	W_stall;
input 	ic_fill_line_5;
input 	i_readdatavalid_d1;
input 	i_readdata_d1_24;
input 	ic_fill_dp_offset_0;
input 	ic_fill_dp_offset_1;
input 	ic_fill_dp_offset_2;
input 	ic_fill_line_0;
input 	ic_fill_line_1;
input 	ic_fill_line_2;
input 	ic_fill_line_3;
input 	ic_fill_line_4;
input 	F_ic_data_rd_addr_nxt_0;
input 	F_ic_data_rd_addr_nxt_1;
input 	F_ic_data_rd_addr_nxt_2;
input 	F_ic_tag_rd_addr_nxt_0;
input 	F_ic_tag_rd_addr_nxt_1;
input 	F_ic_tag_rd_addr_nxt_2;
input 	F_ic_tag_rd_addr_nxt_3;
input 	F_ic_tag_rd_addr_nxt_4;
input 	F_ic_tag_rd_addr_nxt_5;
input 	i_readdata_d1_0;
input 	i_readdata_d1_1;
input 	i_readdata_d1_2;
input 	i_readdata_d1_3;
input 	i_readdata_d1_4;
input 	i_readdata_d1_5;
input 	i_readdata_d1_22;
input 	i_readdata_d1_23;
input 	i_readdata_d1_25;
input 	i_readdata_d1_26;
input 	i_readdata_d1_14;
input 	i_readdata_d1_12;
input 	i_readdata_d1_11;
input 	i_readdata_d1_16;
input 	i_readdata_d1_15;
input 	i_readdata_d1_13;
input 	i_readdata_d1_21;
input 	i_readdata_d1_29;
input 	i_readdata_d1_27;
input 	i_readdata_d1_28;
input 	i_readdata_d1_30;
input 	i_readdata_d1_31;
input 	i_readdata_d1_10;
input 	i_readdata_d1_6;
input 	i_readdata_d1_8;
input 	i_readdata_d1_7;
input 	i_readdata_d1_20;
input 	i_readdata_d1_19;
input 	i_readdata_d1_18;
input 	i_readdata_d1_17;
input 	i_readdata_d1_9;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



processor_altsyncram_1 the_altsyncram(
	.q_b({q_b_31,q_b_30,q_b_29,q_b_28,q_b_27,q_b_26,q_b_25,q_b_24,q_b_23,q_b_22,q_b_21,q_b_20,q_b_19,q_b_18,q_b_17,q_b_16,q_b_15,q_b_14,q_b_13,q_b_12,q_b_11,q_b_10,q_b_9,q_b_8,q_b_7,q_b_6,q_b_5,q_b_4,q_b_3,q_b_2,q_b_1,q_b_0}),
	.rden_b(W_stall),
	.address_a({gnd,gnd,gnd,gnd,ic_fill_line_5,ic_fill_line_4,ic_fill_line_3,ic_fill_line_2,ic_fill_line_1,ic_fill_line_0,ic_fill_dp_offset_2,ic_fill_dp_offset_1,ic_fill_dp_offset_0}),
	.wren_a(i_readdatavalid_d1),
	.data_a({i_readdata_d1_31,i_readdata_d1_30,i_readdata_d1_29,i_readdata_d1_28,i_readdata_d1_27,i_readdata_d1_26,i_readdata_d1_25,i_readdata_d1_24,i_readdata_d1_23,i_readdata_d1_22,i_readdata_d1_21,i_readdata_d1_20,i_readdata_d1_19,i_readdata_d1_18,i_readdata_d1_17,i_readdata_d1_16,
i_readdata_d1_15,i_readdata_d1_14,i_readdata_d1_13,i_readdata_d1_12,i_readdata_d1_11,i_readdata_d1_10,i_readdata_d1_9,i_readdata_d1_8,i_readdata_d1_7,i_readdata_d1_6,i_readdata_d1_5,i_readdata_d1_4,i_readdata_d1_3,i_readdata_d1_2,i_readdata_d1_1,i_readdata_d1_0}),
	.address_b({F_ic_tag_rd_addr_nxt_5,F_ic_tag_rd_addr_nxt_4,F_ic_tag_rd_addr_nxt_3,F_ic_tag_rd_addr_nxt_2,F_ic_tag_rd_addr_nxt_1,F_ic_tag_rd_addr_nxt_0,F_ic_data_rd_addr_nxt_2,F_ic_data_rd_addr_nxt_1,F_ic_data_rd_addr_nxt_0}),
	.clock0(clk_clk));

endmodule

module processor_altsyncram_1 (
	q_b,
	rden_b,
	address_a,
	wren_a,
	data_a,
	address_b,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[31:0] q_b;
input 	rden_b;
input 	[12:0] address_a;
input 	wren_a;
input 	[31:0] data_a;
input 	[8:0] address_b;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



processor_altsyncram_ekj1 auto_generated(
	.q_b({q_b[31],q_b[30],q_b[29],q_b[28],q_b[27],q_b[26],q_b[25],q_b[24],q_b[23],q_b[22],q_b[21],q_b[20],q_b[19],q_b[18],q_b[17],q_b[16],q_b[15],q_b[14],q_b[13],q_b[12],q_b[11],q_b[10],q_b[9],q_b[8],q_b[7],q_b[6],q_b[5],q_b[4],q_b[3],q_b[2],q_b[1],q_b[0]}),
	.rden_b(rden_b),
	.address_a({address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.wren_a(wren_a),
	.data_a({data_a[31],data_a[30],data_a[29],data_a[28],data_a[27],data_a[26],data_a[25],data_a[24],data_a[23],data_a[22],data_a[21],data_a[20],data_a[19],data_a[18],data_a[17],data_a[16],data_a[15],data_a[14],data_a[13],data_a[12],data_a[11],data_a[10],data_a[9],data_a[8],data_a[7],data_a[6],data_a[5],data_a[4],data_a[3],data_a[2],data_a[1],data_a[0]}),
	.address_b({address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.clock0(clock0));

endmodule

module processor_altsyncram_ekj1 (
	q_b,
	rden_b,
	address_a,
	wren_a,
	data_a,
	address_b,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[31:0] q_b;
input 	rden_b;
input 	[8:0] address_a;
input 	wren_a;
input 	[31:0] data_a;
input 	[8:0] address_b;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a24_PORTBDATAOUT_bus;
wire [143:0] ram_block1a0_PORTBDATAOUT_bus;
wire [143:0] ram_block1a1_PORTBDATAOUT_bus;
wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;
wire [143:0] ram_block1a4_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a22_PORTBDATAOUT_bus;
wire [143:0] ram_block1a23_PORTBDATAOUT_bus;
wire [143:0] ram_block1a25_PORTBDATAOUT_bus;
wire [143:0] ram_block1a26_PORTBDATAOUT_bus;
wire [143:0] ram_block1a14_PORTBDATAOUT_bus;
wire [143:0] ram_block1a12_PORTBDATAOUT_bus;
wire [143:0] ram_block1a11_PORTBDATAOUT_bus;
wire [143:0] ram_block1a16_PORTBDATAOUT_bus;
wire [143:0] ram_block1a15_PORTBDATAOUT_bus;
wire [143:0] ram_block1a13_PORTBDATAOUT_bus;
wire [143:0] ram_block1a21_PORTBDATAOUT_bus;
wire [143:0] ram_block1a29_PORTBDATAOUT_bus;
wire [143:0] ram_block1a27_PORTBDATAOUT_bus;
wire [143:0] ram_block1a28_PORTBDATAOUT_bus;
wire [143:0] ram_block1a30_PORTBDATAOUT_bus;
wire [143:0] ram_block1a31_PORTBDATAOUT_bus;
wire [143:0] ram_block1a10_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a8_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a20_PORTBDATAOUT_bus;
wire [143:0] ram_block1a19_PORTBDATAOUT_bus;
wire [143:0] ram_block1a18_PORTBDATAOUT_bus;
wire [143:0] ram_block1a17_PORTBDATAOUT_bus;
wire [143:0] ram_block1a9_PORTBDATAOUT_bus;

assign q_b[24] = ram_block1a24_PORTBDATAOUT_bus[0];

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

assign q_b[2] = ram_block1a2_PORTBDATAOUT_bus[0];

assign q_b[3] = ram_block1a3_PORTBDATAOUT_bus[0];

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[22] = ram_block1a22_PORTBDATAOUT_bus[0];

assign q_b[23] = ram_block1a23_PORTBDATAOUT_bus[0];

assign q_b[25] = ram_block1a25_PORTBDATAOUT_bus[0];

assign q_b[26] = ram_block1a26_PORTBDATAOUT_bus[0];

assign q_b[14] = ram_block1a14_PORTBDATAOUT_bus[0];

assign q_b[12] = ram_block1a12_PORTBDATAOUT_bus[0];

assign q_b[11] = ram_block1a11_PORTBDATAOUT_bus[0];

assign q_b[16] = ram_block1a16_PORTBDATAOUT_bus[0];

assign q_b[15] = ram_block1a15_PORTBDATAOUT_bus[0];

assign q_b[13] = ram_block1a13_PORTBDATAOUT_bus[0];

assign q_b[21] = ram_block1a21_PORTBDATAOUT_bus[0];

assign q_b[29] = ram_block1a29_PORTBDATAOUT_bus[0];

assign q_b[27] = ram_block1a27_PORTBDATAOUT_bus[0];

assign q_b[28] = ram_block1a28_PORTBDATAOUT_bus[0];

assign q_b[30] = ram_block1a30_PORTBDATAOUT_bus[0];

assign q_b[31] = ram_block1a31_PORTBDATAOUT_bus[0];

assign q_b[10] = ram_block1a10_PORTBDATAOUT_bus[0];

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_b[8] = ram_block1a8_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_b[20] = ram_block1a20_PORTBDATAOUT_bus[0];

assign q_b[19] = ram_block1a19_PORTBDATAOUT_bus[0];

assign q_b[18] = ram_block1a18_PORTBDATAOUT_bus[0];

assign q_b[17] = ram_block1a17_PORTBDATAOUT_bus[0];

assign q_b[9] = ram_block1a9_PORTBDATAOUT_bus[0];

cyclonev_ram_block ram_block1a24(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(rden_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[24]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a24_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a24.clk0_core_clock_enable = "ena0";
defparam ram_block1a24.clk1_core_clock_enable = "ena1";
defparam ram_block1a24.data_interleave_offset_in_bits = 1;
defparam ram_block1a24.data_interleave_width_in_bits = 1;
defparam ram_block1a24.logical_ram_name = "processor_cpu:cpu|processor_cpu_ic_data_module:processor_cpu_ic_data|altsyncram:the_altsyncram|altsyncram_ekj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a24.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a24.operation_mode = "dual_port";
defparam ram_block1a24.port_a_address_clear = "none";
defparam ram_block1a24.port_a_address_width = 9;
defparam ram_block1a24.port_a_data_out_clear = "none";
defparam ram_block1a24.port_a_data_out_clock = "none";
defparam ram_block1a24.port_a_data_width = 1;
defparam ram_block1a24.port_a_first_address = 0;
defparam ram_block1a24.port_a_first_bit_number = 24;
defparam ram_block1a24.port_a_last_address = 511;
defparam ram_block1a24.port_a_logical_ram_depth = 512;
defparam ram_block1a24.port_a_logical_ram_width = 32;
defparam ram_block1a24.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a24.port_b_address_clear = "none";
defparam ram_block1a24.port_b_address_clock = "clock1";
defparam ram_block1a24.port_b_address_width = 9;
defparam ram_block1a24.port_b_data_out_clear = "none";
defparam ram_block1a24.port_b_data_out_clock = "none";
defparam ram_block1a24.port_b_data_width = 1;
defparam ram_block1a24.port_b_first_address = 0;
defparam ram_block1a24.port_b_first_bit_number = 24;
defparam ram_block1a24.port_b_last_address = 511;
defparam ram_block1a24.port_b_logical_ram_depth = 512;
defparam ram_block1a24.port_b_logical_ram_width = 32;
defparam ram_block1a24.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a24.port_b_read_enable_clock = "clock1";
defparam ram_block1a24.ram_block_type = "auto";

cyclonev_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(rden_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.clk1_core_clock_enable = "ena1";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.logical_ram_name = "processor_cpu:cpu|processor_cpu_ic_data_module:processor_cpu_ic_data|altsyncram:the_altsyncram|altsyncram_ekj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a0.operation_mode = "dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 9;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 511;
defparam ram_block1a0.port_a_logical_ram_depth = 512;
defparam ram_block1a0.port_a_logical_ram_width = 32;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_address_clear = "none";
defparam ram_block1a0.port_b_address_clock = "clock1";
defparam ram_block1a0.port_b_address_width = 9;
defparam ram_block1a0.port_b_data_out_clear = "none";
defparam ram_block1a0.port_b_data_out_clock = "none";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 511;
defparam ram_block1a0.port_b_logical_ram_depth = 512;
defparam ram_block1a0.port_b_logical_ram_width = 32;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock1";
defparam ram_block1a0.ram_block_type = "auto";

cyclonev_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(rden_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a1.clk0_core_clock_enable = "ena0";
defparam ram_block1a1.clk1_core_clock_enable = "ena1";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.logical_ram_name = "processor_cpu:cpu|processor_cpu_ic_data_module:processor_cpu_ic_data|altsyncram:the_altsyncram|altsyncram_ekj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a1.operation_mode = "dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 9;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 511;
defparam ram_block1a1.port_a_logical_ram_depth = 512;
defparam ram_block1a1.port_a_logical_ram_width = 32;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_address_clear = "none";
defparam ram_block1a1.port_b_address_clock = "clock1";
defparam ram_block1a1.port_b_address_width = 9;
defparam ram_block1a1.port_b_data_out_clear = "none";
defparam ram_block1a1.port_b_data_out_clock = "none";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 511;
defparam ram_block1a1.port_b_logical_ram_depth = 512;
defparam ram_block1a1.port_b_logical_ram_width = 32;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock1";
defparam ram_block1a1.ram_block_type = "auto";

cyclonev_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(rden_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a2.clk0_core_clock_enable = "ena0";
defparam ram_block1a2.clk1_core_clock_enable = "ena1";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.logical_ram_name = "processor_cpu:cpu|processor_cpu_ic_data_module:processor_cpu_ic_data|altsyncram:the_altsyncram|altsyncram_ekj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a2.operation_mode = "dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 9;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 511;
defparam ram_block1a2.port_a_logical_ram_depth = 512;
defparam ram_block1a2.port_a_logical_ram_width = 32;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_address_clear = "none";
defparam ram_block1a2.port_b_address_clock = "clock1";
defparam ram_block1a2.port_b_address_width = 9;
defparam ram_block1a2.port_b_data_out_clear = "none";
defparam ram_block1a2.port_b_data_out_clock = "none";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 511;
defparam ram_block1a2.port_b_logical_ram_depth = 512;
defparam ram_block1a2.port_b_logical_ram_width = 32;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock1";
defparam ram_block1a2.ram_block_type = "auto";

cyclonev_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(rden_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a3.clk0_core_clock_enable = "ena0";
defparam ram_block1a3.clk1_core_clock_enable = "ena1";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.logical_ram_name = "processor_cpu:cpu|processor_cpu_ic_data_module:processor_cpu_ic_data|altsyncram:the_altsyncram|altsyncram_ekj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a3.operation_mode = "dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 9;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 511;
defparam ram_block1a3.port_a_logical_ram_depth = 512;
defparam ram_block1a3.port_a_logical_ram_width = 32;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_address_clear = "none";
defparam ram_block1a3.port_b_address_clock = "clock1";
defparam ram_block1a3.port_b_address_width = 9;
defparam ram_block1a3.port_b_data_out_clear = "none";
defparam ram_block1a3.port_b_data_out_clock = "none";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 511;
defparam ram_block1a3.port_b_logical_ram_depth = 512;
defparam ram_block1a3.port_b_logical_ram_width = 32;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock1";
defparam ram_block1a3.ram_block_type = "auto";

cyclonev_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(rden_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a4.clk0_core_clock_enable = "ena0";
defparam ram_block1a4.clk1_core_clock_enable = "ena1";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.logical_ram_name = "processor_cpu:cpu|processor_cpu_ic_data_module:processor_cpu_ic_data|altsyncram:the_altsyncram|altsyncram_ekj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a4.operation_mode = "dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 9;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 511;
defparam ram_block1a4.port_a_logical_ram_depth = 512;
defparam ram_block1a4.port_a_logical_ram_width = 32;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_address_clear = "none";
defparam ram_block1a4.port_b_address_clock = "clock1";
defparam ram_block1a4.port_b_address_width = 9;
defparam ram_block1a4.port_b_data_out_clear = "none";
defparam ram_block1a4.port_b_data_out_clock = "none";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 511;
defparam ram_block1a4.port_b_logical_ram_depth = 512;
defparam ram_block1a4.port_b_logical_ram_width = 32;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock1";
defparam ram_block1a4.ram_block_type = "auto";

cyclonev_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(rden_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a5.clk0_core_clock_enable = "ena0";
defparam ram_block1a5.clk1_core_clock_enable = "ena1";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "processor_cpu:cpu|processor_cpu_ic_data_module:processor_cpu_ic_data|altsyncram:the_altsyncram|altsyncram_ekj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 9;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 511;
defparam ram_block1a5.port_a_logical_ram_depth = 512;
defparam ram_block1a5.port_a_logical_ram_width = 32;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_address_clear = "none";
defparam ram_block1a5.port_b_address_clock = "clock1";
defparam ram_block1a5.port_b_address_width = 9;
defparam ram_block1a5.port_b_data_out_clear = "none";
defparam ram_block1a5.port_b_data_out_clock = "none";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 511;
defparam ram_block1a5.port_b_logical_ram_depth = 512;
defparam ram_block1a5.port_b_logical_ram_width = 32;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock1";
defparam ram_block1a5.ram_block_type = "auto";

cyclonev_ram_block ram_block1a22(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(rden_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[22]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a22_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a22.clk0_core_clock_enable = "ena0";
defparam ram_block1a22.clk1_core_clock_enable = "ena1";
defparam ram_block1a22.data_interleave_offset_in_bits = 1;
defparam ram_block1a22.data_interleave_width_in_bits = 1;
defparam ram_block1a22.logical_ram_name = "processor_cpu:cpu|processor_cpu_ic_data_module:processor_cpu_ic_data|altsyncram:the_altsyncram|altsyncram_ekj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a22.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a22.operation_mode = "dual_port";
defparam ram_block1a22.port_a_address_clear = "none";
defparam ram_block1a22.port_a_address_width = 9;
defparam ram_block1a22.port_a_data_out_clear = "none";
defparam ram_block1a22.port_a_data_out_clock = "none";
defparam ram_block1a22.port_a_data_width = 1;
defparam ram_block1a22.port_a_first_address = 0;
defparam ram_block1a22.port_a_first_bit_number = 22;
defparam ram_block1a22.port_a_last_address = 511;
defparam ram_block1a22.port_a_logical_ram_depth = 512;
defparam ram_block1a22.port_a_logical_ram_width = 32;
defparam ram_block1a22.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a22.port_b_address_clear = "none";
defparam ram_block1a22.port_b_address_clock = "clock1";
defparam ram_block1a22.port_b_address_width = 9;
defparam ram_block1a22.port_b_data_out_clear = "none";
defparam ram_block1a22.port_b_data_out_clock = "none";
defparam ram_block1a22.port_b_data_width = 1;
defparam ram_block1a22.port_b_first_address = 0;
defparam ram_block1a22.port_b_first_bit_number = 22;
defparam ram_block1a22.port_b_last_address = 511;
defparam ram_block1a22.port_b_logical_ram_depth = 512;
defparam ram_block1a22.port_b_logical_ram_width = 32;
defparam ram_block1a22.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a22.port_b_read_enable_clock = "clock1";
defparam ram_block1a22.ram_block_type = "auto";

cyclonev_ram_block ram_block1a23(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(rden_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[23]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a23_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a23.clk0_core_clock_enable = "ena0";
defparam ram_block1a23.clk1_core_clock_enable = "ena1";
defparam ram_block1a23.data_interleave_offset_in_bits = 1;
defparam ram_block1a23.data_interleave_width_in_bits = 1;
defparam ram_block1a23.logical_ram_name = "processor_cpu:cpu|processor_cpu_ic_data_module:processor_cpu_ic_data|altsyncram:the_altsyncram|altsyncram_ekj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a23.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a23.operation_mode = "dual_port";
defparam ram_block1a23.port_a_address_clear = "none";
defparam ram_block1a23.port_a_address_width = 9;
defparam ram_block1a23.port_a_data_out_clear = "none";
defparam ram_block1a23.port_a_data_out_clock = "none";
defparam ram_block1a23.port_a_data_width = 1;
defparam ram_block1a23.port_a_first_address = 0;
defparam ram_block1a23.port_a_first_bit_number = 23;
defparam ram_block1a23.port_a_last_address = 511;
defparam ram_block1a23.port_a_logical_ram_depth = 512;
defparam ram_block1a23.port_a_logical_ram_width = 32;
defparam ram_block1a23.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a23.port_b_address_clear = "none";
defparam ram_block1a23.port_b_address_clock = "clock1";
defparam ram_block1a23.port_b_address_width = 9;
defparam ram_block1a23.port_b_data_out_clear = "none";
defparam ram_block1a23.port_b_data_out_clock = "none";
defparam ram_block1a23.port_b_data_width = 1;
defparam ram_block1a23.port_b_first_address = 0;
defparam ram_block1a23.port_b_first_bit_number = 23;
defparam ram_block1a23.port_b_last_address = 511;
defparam ram_block1a23.port_b_logical_ram_depth = 512;
defparam ram_block1a23.port_b_logical_ram_width = 32;
defparam ram_block1a23.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a23.port_b_read_enable_clock = "clock1";
defparam ram_block1a23.ram_block_type = "auto";

cyclonev_ram_block ram_block1a25(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(rden_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[25]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a25_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a25.clk0_core_clock_enable = "ena0";
defparam ram_block1a25.clk1_core_clock_enable = "ena1";
defparam ram_block1a25.data_interleave_offset_in_bits = 1;
defparam ram_block1a25.data_interleave_width_in_bits = 1;
defparam ram_block1a25.logical_ram_name = "processor_cpu:cpu|processor_cpu_ic_data_module:processor_cpu_ic_data|altsyncram:the_altsyncram|altsyncram_ekj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a25.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a25.operation_mode = "dual_port";
defparam ram_block1a25.port_a_address_clear = "none";
defparam ram_block1a25.port_a_address_width = 9;
defparam ram_block1a25.port_a_data_out_clear = "none";
defparam ram_block1a25.port_a_data_out_clock = "none";
defparam ram_block1a25.port_a_data_width = 1;
defparam ram_block1a25.port_a_first_address = 0;
defparam ram_block1a25.port_a_first_bit_number = 25;
defparam ram_block1a25.port_a_last_address = 511;
defparam ram_block1a25.port_a_logical_ram_depth = 512;
defparam ram_block1a25.port_a_logical_ram_width = 32;
defparam ram_block1a25.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a25.port_b_address_clear = "none";
defparam ram_block1a25.port_b_address_clock = "clock1";
defparam ram_block1a25.port_b_address_width = 9;
defparam ram_block1a25.port_b_data_out_clear = "none";
defparam ram_block1a25.port_b_data_out_clock = "none";
defparam ram_block1a25.port_b_data_width = 1;
defparam ram_block1a25.port_b_first_address = 0;
defparam ram_block1a25.port_b_first_bit_number = 25;
defparam ram_block1a25.port_b_last_address = 511;
defparam ram_block1a25.port_b_logical_ram_depth = 512;
defparam ram_block1a25.port_b_logical_ram_width = 32;
defparam ram_block1a25.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a25.port_b_read_enable_clock = "clock1";
defparam ram_block1a25.ram_block_type = "auto";

cyclonev_ram_block ram_block1a26(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(rden_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[26]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a26_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a26.clk0_core_clock_enable = "ena0";
defparam ram_block1a26.clk1_core_clock_enable = "ena1";
defparam ram_block1a26.data_interleave_offset_in_bits = 1;
defparam ram_block1a26.data_interleave_width_in_bits = 1;
defparam ram_block1a26.logical_ram_name = "processor_cpu:cpu|processor_cpu_ic_data_module:processor_cpu_ic_data|altsyncram:the_altsyncram|altsyncram_ekj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a26.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a26.operation_mode = "dual_port";
defparam ram_block1a26.port_a_address_clear = "none";
defparam ram_block1a26.port_a_address_width = 9;
defparam ram_block1a26.port_a_data_out_clear = "none";
defparam ram_block1a26.port_a_data_out_clock = "none";
defparam ram_block1a26.port_a_data_width = 1;
defparam ram_block1a26.port_a_first_address = 0;
defparam ram_block1a26.port_a_first_bit_number = 26;
defparam ram_block1a26.port_a_last_address = 511;
defparam ram_block1a26.port_a_logical_ram_depth = 512;
defparam ram_block1a26.port_a_logical_ram_width = 32;
defparam ram_block1a26.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a26.port_b_address_clear = "none";
defparam ram_block1a26.port_b_address_clock = "clock1";
defparam ram_block1a26.port_b_address_width = 9;
defparam ram_block1a26.port_b_data_out_clear = "none";
defparam ram_block1a26.port_b_data_out_clock = "none";
defparam ram_block1a26.port_b_data_width = 1;
defparam ram_block1a26.port_b_first_address = 0;
defparam ram_block1a26.port_b_first_bit_number = 26;
defparam ram_block1a26.port_b_last_address = 511;
defparam ram_block1a26.port_b_logical_ram_depth = 512;
defparam ram_block1a26.port_b_logical_ram_width = 32;
defparam ram_block1a26.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a26.port_b_read_enable_clock = "clock1";
defparam ram_block1a26.ram_block_type = "auto";

cyclonev_ram_block ram_block1a14(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(rden_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a14_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a14.clk0_core_clock_enable = "ena0";
defparam ram_block1a14.clk1_core_clock_enable = "ena1";
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.logical_ram_name = "processor_cpu:cpu|processor_cpu_ic_data_module:processor_cpu_ic_data|altsyncram:the_altsyncram|altsyncram_ekj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a14.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a14.operation_mode = "dual_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 9;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 511;
defparam ram_block1a14.port_a_logical_ram_depth = 512;
defparam ram_block1a14.port_a_logical_ram_width = 32;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a14.port_b_address_clear = "none";
defparam ram_block1a14.port_b_address_clock = "clock1";
defparam ram_block1a14.port_b_address_width = 9;
defparam ram_block1a14.port_b_data_out_clear = "none";
defparam ram_block1a14.port_b_data_out_clock = "none";
defparam ram_block1a14.port_b_data_width = 1;
defparam ram_block1a14.port_b_first_address = 0;
defparam ram_block1a14.port_b_first_bit_number = 14;
defparam ram_block1a14.port_b_last_address = 511;
defparam ram_block1a14.port_b_logical_ram_depth = 512;
defparam ram_block1a14.port_b_logical_ram_width = 32;
defparam ram_block1a14.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a14.port_b_read_enable_clock = "clock1";
defparam ram_block1a14.ram_block_type = "auto";

cyclonev_ram_block ram_block1a12(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(rden_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a12_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a12.clk0_core_clock_enable = "ena0";
defparam ram_block1a12.clk1_core_clock_enable = "ena1";
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.logical_ram_name = "processor_cpu:cpu|processor_cpu_ic_data_module:processor_cpu_ic_data|altsyncram:the_altsyncram|altsyncram_ekj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a12.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a12.operation_mode = "dual_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 9;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 511;
defparam ram_block1a12.port_a_logical_ram_depth = 512;
defparam ram_block1a12.port_a_logical_ram_width = 32;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a12.port_b_address_clear = "none";
defparam ram_block1a12.port_b_address_clock = "clock1";
defparam ram_block1a12.port_b_address_width = 9;
defparam ram_block1a12.port_b_data_out_clear = "none";
defparam ram_block1a12.port_b_data_out_clock = "none";
defparam ram_block1a12.port_b_data_width = 1;
defparam ram_block1a12.port_b_first_address = 0;
defparam ram_block1a12.port_b_first_bit_number = 12;
defparam ram_block1a12.port_b_last_address = 511;
defparam ram_block1a12.port_b_logical_ram_depth = 512;
defparam ram_block1a12.port_b_logical_ram_width = 32;
defparam ram_block1a12.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a12.port_b_read_enable_clock = "clock1";
defparam ram_block1a12.ram_block_type = "auto";

cyclonev_ram_block ram_block1a11(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(rden_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a11_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a11.clk0_core_clock_enable = "ena0";
defparam ram_block1a11.clk1_core_clock_enable = "ena1";
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.logical_ram_name = "processor_cpu:cpu|processor_cpu_ic_data_module:processor_cpu_ic_data|altsyncram:the_altsyncram|altsyncram_ekj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a11.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a11.operation_mode = "dual_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 9;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 511;
defparam ram_block1a11.port_a_logical_ram_depth = 512;
defparam ram_block1a11.port_a_logical_ram_width = 32;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a11.port_b_address_clear = "none";
defparam ram_block1a11.port_b_address_clock = "clock1";
defparam ram_block1a11.port_b_address_width = 9;
defparam ram_block1a11.port_b_data_out_clear = "none";
defparam ram_block1a11.port_b_data_out_clock = "none";
defparam ram_block1a11.port_b_data_width = 1;
defparam ram_block1a11.port_b_first_address = 0;
defparam ram_block1a11.port_b_first_bit_number = 11;
defparam ram_block1a11.port_b_last_address = 511;
defparam ram_block1a11.port_b_logical_ram_depth = 512;
defparam ram_block1a11.port_b_logical_ram_width = 32;
defparam ram_block1a11.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a11.port_b_read_enable_clock = "clock1";
defparam ram_block1a11.ram_block_type = "auto";

cyclonev_ram_block ram_block1a16(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(rden_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a16_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a16.clk0_core_clock_enable = "ena0";
defparam ram_block1a16.clk1_core_clock_enable = "ena1";
defparam ram_block1a16.data_interleave_offset_in_bits = 1;
defparam ram_block1a16.data_interleave_width_in_bits = 1;
defparam ram_block1a16.logical_ram_name = "processor_cpu:cpu|processor_cpu_ic_data_module:processor_cpu_ic_data|altsyncram:the_altsyncram|altsyncram_ekj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a16.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a16.operation_mode = "dual_port";
defparam ram_block1a16.port_a_address_clear = "none";
defparam ram_block1a16.port_a_address_width = 9;
defparam ram_block1a16.port_a_data_out_clear = "none";
defparam ram_block1a16.port_a_data_out_clock = "none";
defparam ram_block1a16.port_a_data_width = 1;
defparam ram_block1a16.port_a_first_address = 0;
defparam ram_block1a16.port_a_first_bit_number = 16;
defparam ram_block1a16.port_a_last_address = 511;
defparam ram_block1a16.port_a_logical_ram_depth = 512;
defparam ram_block1a16.port_a_logical_ram_width = 32;
defparam ram_block1a16.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a16.port_b_address_clear = "none";
defparam ram_block1a16.port_b_address_clock = "clock1";
defparam ram_block1a16.port_b_address_width = 9;
defparam ram_block1a16.port_b_data_out_clear = "none";
defparam ram_block1a16.port_b_data_out_clock = "none";
defparam ram_block1a16.port_b_data_width = 1;
defparam ram_block1a16.port_b_first_address = 0;
defparam ram_block1a16.port_b_first_bit_number = 16;
defparam ram_block1a16.port_b_last_address = 511;
defparam ram_block1a16.port_b_logical_ram_depth = 512;
defparam ram_block1a16.port_b_logical_ram_width = 32;
defparam ram_block1a16.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a16.port_b_read_enable_clock = "clock1";
defparam ram_block1a16.ram_block_type = "auto";

cyclonev_ram_block ram_block1a15(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(rden_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a15_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a15.clk0_core_clock_enable = "ena0";
defparam ram_block1a15.clk1_core_clock_enable = "ena1";
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.logical_ram_name = "processor_cpu:cpu|processor_cpu_ic_data_module:processor_cpu_ic_data|altsyncram:the_altsyncram|altsyncram_ekj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a15.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a15.operation_mode = "dual_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 9;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 511;
defparam ram_block1a15.port_a_logical_ram_depth = 512;
defparam ram_block1a15.port_a_logical_ram_width = 32;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a15.port_b_address_clear = "none";
defparam ram_block1a15.port_b_address_clock = "clock1";
defparam ram_block1a15.port_b_address_width = 9;
defparam ram_block1a15.port_b_data_out_clear = "none";
defparam ram_block1a15.port_b_data_out_clock = "none";
defparam ram_block1a15.port_b_data_width = 1;
defparam ram_block1a15.port_b_first_address = 0;
defparam ram_block1a15.port_b_first_bit_number = 15;
defparam ram_block1a15.port_b_last_address = 511;
defparam ram_block1a15.port_b_logical_ram_depth = 512;
defparam ram_block1a15.port_b_logical_ram_width = 32;
defparam ram_block1a15.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a15.port_b_read_enable_clock = "clock1";
defparam ram_block1a15.ram_block_type = "auto";

cyclonev_ram_block ram_block1a13(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(rden_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a13_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a13.clk0_core_clock_enable = "ena0";
defparam ram_block1a13.clk1_core_clock_enable = "ena1";
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.logical_ram_name = "processor_cpu:cpu|processor_cpu_ic_data_module:processor_cpu_ic_data|altsyncram:the_altsyncram|altsyncram_ekj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a13.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a13.operation_mode = "dual_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 9;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 511;
defparam ram_block1a13.port_a_logical_ram_depth = 512;
defparam ram_block1a13.port_a_logical_ram_width = 32;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a13.port_b_address_clear = "none";
defparam ram_block1a13.port_b_address_clock = "clock1";
defparam ram_block1a13.port_b_address_width = 9;
defparam ram_block1a13.port_b_data_out_clear = "none";
defparam ram_block1a13.port_b_data_out_clock = "none";
defparam ram_block1a13.port_b_data_width = 1;
defparam ram_block1a13.port_b_first_address = 0;
defparam ram_block1a13.port_b_first_bit_number = 13;
defparam ram_block1a13.port_b_last_address = 511;
defparam ram_block1a13.port_b_logical_ram_depth = 512;
defparam ram_block1a13.port_b_logical_ram_width = 32;
defparam ram_block1a13.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a13.port_b_read_enable_clock = "clock1";
defparam ram_block1a13.ram_block_type = "auto";

cyclonev_ram_block ram_block1a21(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(rden_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[21]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a21_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a21.clk0_core_clock_enable = "ena0";
defparam ram_block1a21.clk1_core_clock_enable = "ena1";
defparam ram_block1a21.data_interleave_offset_in_bits = 1;
defparam ram_block1a21.data_interleave_width_in_bits = 1;
defparam ram_block1a21.logical_ram_name = "processor_cpu:cpu|processor_cpu_ic_data_module:processor_cpu_ic_data|altsyncram:the_altsyncram|altsyncram_ekj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a21.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a21.operation_mode = "dual_port";
defparam ram_block1a21.port_a_address_clear = "none";
defparam ram_block1a21.port_a_address_width = 9;
defparam ram_block1a21.port_a_data_out_clear = "none";
defparam ram_block1a21.port_a_data_out_clock = "none";
defparam ram_block1a21.port_a_data_width = 1;
defparam ram_block1a21.port_a_first_address = 0;
defparam ram_block1a21.port_a_first_bit_number = 21;
defparam ram_block1a21.port_a_last_address = 511;
defparam ram_block1a21.port_a_logical_ram_depth = 512;
defparam ram_block1a21.port_a_logical_ram_width = 32;
defparam ram_block1a21.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a21.port_b_address_clear = "none";
defparam ram_block1a21.port_b_address_clock = "clock1";
defparam ram_block1a21.port_b_address_width = 9;
defparam ram_block1a21.port_b_data_out_clear = "none";
defparam ram_block1a21.port_b_data_out_clock = "none";
defparam ram_block1a21.port_b_data_width = 1;
defparam ram_block1a21.port_b_first_address = 0;
defparam ram_block1a21.port_b_first_bit_number = 21;
defparam ram_block1a21.port_b_last_address = 511;
defparam ram_block1a21.port_b_logical_ram_depth = 512;
defparam ram_block1a21.port_b_logical_ram_width = 32;
defparam ram_block1a21.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a21.port_b_read_enable_clock = "clock1";
defparam ram_block1a21.ram_block_type = "auto";

cyclonev_ram_block ram_block1a29(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(rden_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[29]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a29_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a29.clk0_core_clock_enable = "ena0";
defparam ram_block1a29.clk1_core_clock_enable = "ena1";
defparam ram_block1a29.data_interleave_offset_in_bits = 1;
defparam ram_block1a29.data_interleave_width_in_bits = 1;
defparam ram_block1a29.logical_ram_name = "processor_cpu:cpu|processor_cpu_ic_data_module:processor_cpu_ic_data|altsyncram:the_altsyncram|altsyncram_ekj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a29.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a29.operation_mode = "dual_port";
defparam ram_block1a29.port_a_address_clear = "none";
defparam ram_block1a29.port_a_address_width = 9;
defparam ram_block1a29.port_a_data_out_clear = "none";
defparam ram_block1a29.port_a_data_out_clock = "none";
defparam ram_block1a29.port_a_data_width = 1;
defparam ram_block1a29.port_a_first_address = 0;
defparam ram_block1a29.port_a_first_bit_number = 29;
defparam ram_block1a29.port_a_last_address = 511;
defparam ram_block1a29.port_a_logical_ram_depth = 512;
defparam ram_block1a29.port_a_logical_ram_width = 32;
defparam ram_block1a29.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a29.port_b_address_clear = "none";
defparam ram_block1a29.port_b_address_clock = "clock1";
defparam ram_block1a29.port_b_address_width = 9;
defparam ram_block1a29.port_b_data_out_clear = "none";
defparam ram_block1a29.port_b_data_out_clock = "none";
defparam ram_block1a29.port_b_data_width = 1;
defparam ram_block1a29.port_b_first_address = 0;
defparam ram_block1a29.port_b_first_bit_number = 29;
defparam ram_block1a29.port_b_last_address = 511;
defparam ram_block1a29.port_b_logical_ram_depth = 512;
defparam ram_block1a29.port_b_logical_ram_width = 32;
defparam ram_block1a29.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a29.port_b_read_enable_clock = "clock1";
defparam ram_block1a29.ram_block_type = "auto";

cyclonev_ram_block ram_block1a27(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(rden_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[27]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a27_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a27.clk0_core_clock_enable = "ena0";
defparam ram_block1a27.clk1_core_clock_enable = "ena1";
defparam ram_block1a27.data_interleave_offset_in_bits = 1;
defparam ram_block1a27.data_interleave_width_in_bits = 1;
defparam ram_block1a27.logical_ram_name = "processor_cpu:cpu|processor_cpu_ic_data_module:processor_cpu_ic_data|altsyncram:the_altsyncram|altsyncram_ekj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a27.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a27.operation_mode = "dual_port";
defparam ram_block1a27.port_a_address_clear = "none";
defparam ram_block1a27.port_a_address_width = 9;
defparam ram_block1a27.port_a_data_out_clear = "none";
defparam ram_block1a27.port_a_data_out_clock = "none";
defparam ram_block1a27.port_a_data_width = 1;
defparam ram_block1a27.port_a_first_address = 0;
defparam ram_block1a27.port_a_first_bit_number = 27;
defparam ram_block1a27.port_a_last_address = 511;
defparam ram_block1a27.port_a_logical_ram_depth = 512;
defparam ram_block1a27.port_a_logical_ram_width = 32;
defparam ram_block1a27.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a27.port_b_address_clear = "none";
defparam ram_block1a27.port_b_address_clock = "clock1";
defparam ram_block1a27.port_b_address_width = 9;
defparam ram_block1a27.port_b_data_out_clear = "none";
defparam ram_block1a27.port_b_data_out_clock = "none";
defparam ram_block1a27.port_b_data_width = 1;
defparam ram_block1a27.port_b_first_address = 0;
defparam ram_block1a27.port_b_first_bit_number = 27;
defparam ram_block1a27.port_b_last_address = 511;
defparam ram_block1a27.port_b_logical_ram_depth = 512;
defparam ram_block1a27.port_b_logical_ram_width = 32;
defparam ram_block1a27.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a27.port_b_read_enable_clock = "clock1";
defparam ram_block1a27.ram_block_type = "auto";

cyclonev_ram_block ram_block1a28(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(rden_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[28]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a28_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a28.clk0_core_clock_enable = "ena0";
defparam ram_block1a28.clk1_core_clock_enable = "ena1";
defparam ram_block1a28.data_interleave_offset_in_bits = 1;
defparam ram_block1a28.data_interleave_width_in_bits = 1;
defparam ram_block1a28.logical_ram_name = "processor_cpu:cpu|processor_cpu_ic_data_module:processor_cpu_ic_data|altsyncram:the_altsyncram|altsyncram_ekj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a28.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a28.operation_mode = "dual_port";
defparam ram_block1a28.port_a_address_clear = "none";
defparam ram_block1a28.port_a_address_width = 9;
defparam ram_block1a28.port_a_data_out_clear = "none";
defparam ram_block1a28.port_a_data_out_clock = "none";
defparam ram_block1a28.port_a_data_width = 1;
defparam ram_block1a28.port_a_first_address = 0;
defparam ram_block1a28.port_a_first_bit_number = 28;
defparam ram_block1a28.port_a_last_address = 511;
defparam ram_block1a28.port_a_logical_ram_depth = 512;
defparam ram_block1a28.port_a_logical_ram_width = 32;
defparam ram_block1a28.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a28.port_b_address_clear = "none";
defparam ram_block1a28.port_b_address_clock = "clock1";
defparam ram_block1a28.port_b_address_width = 9;
defparam ram_block1a28.port_b_data_out_clear = "none";
defparam ram_block1a28.port_b_data_out_clock = "none";
defparam ram_block1a28.port_b_data_width = 1;
defparam ram_block1a28.port_b_first_address = 0;
defparam ram_block1a28.port_b_first_bit_number = 28;
defparam ram_block1a28.port_b_last_address = 511;
defparam ram_block1a28.port_b_logical_ram_depth = 512;
defparam ram_block1a28.port_b_logical_ram_width = 32;
defparam ram_block1a28.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a28.port_b_read_enable_clock = "clock1";
defparam ram_block1a28.ram_block_type = "auto";

cyclonev_ram_block ram_block1a30(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(rden_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[30]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a30_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a30.clk0_core_clock_enable = "ena0";
defparam ram_block1a30.clk1_core_clock_enable = "ena1";
defparam ram_block1a30.data_interleave_offset_in_bits = 1;
defparam ram_block1a30.data_interleave_width_in_bits = 1;
defparam ram_block1a30.logical_ram_name = "processor_cpu:cpu|processor_cpu_ic_data_module:processor_cpu_ic_data|altsyncram:the_altsyncram|altsyncram_ekj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a30.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a30.operation_mode = "dual_port";
defparam ram_block1a30.port_a_address_clear = "none";
defparam ram_block1a30.port_a_address_width = 9;
defparam ram_block1a30.port_a_data_out_clear = "none";
defparam ram_block1a30.port_a_data_out_clock = "none";
defparam ram_block1a30.port_a_data_width = 1;
defparam ram_block1a30.port_a_first_address = 0;
defparam ram_block1a30.port_a_first_bit_number = 30;
defparam ram_block1a30.port_a_last_address = 511;
defparam ram_block1a30.port_a_logical_ram_depth = 512;
defparam ram_block1a30.port_a_logical_ram_width = 32;
defparam ram_block1a30.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a30.port_b_address_clear = "none";
defparam ram_block1a30.port_b_address_clock = "clock1";
defparam ram_block1a30.port_b_address_width = 9;
defparam ram_block1a30.port_b_data_out_clear = "none";
defparam ram_block1a30.port_b_data_out_clock = "none";
defparam ram_block1a30.port_b_data_width = 1;
defparam ram_block1a30.port_b_first_address = 0;
defparam ram_block1a30.port_b_first_bit_number = 30;
defparam ram_block1a30.port_b_last_address = 511;
defparam ram_block1a30.port_b_logical_ram_depth = 512;
defparam ram_block1a30.port_b_logical_ram_width = 32;
defparam ram_block1a30.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a30.port_b_read_enable_clock = "clock1";
defparam ram_block1a30.ram_block_type = "auto";

cyclonev_ram_block ram_block1a31(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(rden_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[31]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a31_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a31.clk0_core_clock_enable = "ena0";
defparam ram_block1a31.clk1_core_clock_enable = "ena1";
defparam ram_block1a31.data_interleave_offset_in_bits = 1;
defparam ram_block1a31.data_interleave_width_in_bits = 1;
defparam ram_block1a31.logical_ram_name = "processor_cpu:cpu|processor_cpu_ic_data_module:processor_cpu_ic_data|altsyncram:the_altsyncram|altsyncram_ekj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a31.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a31.operation_mode = "dual_port";
defparam ram_block1a31.port_a_address_clear = "none";
defparam ram_block1a31.port_a_address_width = 9;
defparam ram_block1a31.port_a_data_out_clear = "none";
defparam ram_block1a31.port_a_data_out_clock = "none";
defparam ram_block1a31.port_a_data_width = 1;
defparam ram_block1a31.port_a_first_address = 0;
defparam ram_block1a31.port_a_first_bit_number = 31;
defparam ram_block1a31.port_a_last_address = 511;
defparam ram_block1a31.port_a_logical_ram_depth = 512;
defparam ram_block1a31.port_a_logical_ram_width = 32;
defparam ram_block1a31.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a31.port_b_address_clear = "none";
defparam ram_block1a31.port_b_address_clock = "clock1";
defparam ram_block1a31.port_b_address_width = 9;
defparam ram_block1a31.port_b_data_out_clear = "none";
defparam ram_block1a31.port_b_data_out_clock = "none";
defparam ram_block1a31.port_b_data_width = 1;
defparam ram_block1a31.port_b_first_address = 0;
defparam ram_block1a31.port_b_first_bit_number = 31;
defparam ram_block1a31.port_b_last_address = 511;
defparam ram_block1a31.port_b_logical_ram_depth = 512;
defparam ram_block1a31.port_b_logical_ram_width = 32;
defparam ram_block1a31.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a31.port_b_read_enable_clock = "clock1";
defparam ram_block1a31.ram_block_type = "auto";

cyclonev_ram_block ram_block1a10(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(rden_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a10_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a10.clk0_core_clock_enable = "ena0";
defparam ram_block1a10.clk1_core_clock_enable = "ena1";
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.logical_ram_name = "processor_cpu:cpu|processor_cpu_ic_data_module:processor_cpu_ic_data|altsyncram:the_altsyncram|altsyncram_ekj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a10.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a10.operation_mode = "dual_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 9;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 511;
defparam ram_block1a10.port_a_logical_ram_depth = 512;
defparam ram_block1a10.port_a_logical_ram_width = 32;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a10.port_b_address_clear = "none";
defparam ram_block1a10.port_b_address_clock = "clock1";
defparam ram_block1a10.port_b_address_width = 9;
defparam ram_block1a10.port_b_data_out_clear = "none";
defparam ram_block1a10.port_b_data_out_clock = "none";
defparam ram_block1a10.port_b_data_width = 1;
defparam ram_block1a10.port_b_first_address = 0;
defparam ram_block1a10.port_b_first_bit_number = 10;
defparam ram_block1a10.port_b_last_address = 511;
defparam ram_block1a10.port_b_logical_ram_depth = 512;
defparam ram_block1a10.port_b_logical_ram_width = 32;
defparam ram_block1a10.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a10.port_b_read_enable_clock = "clock1";
defparam ram_block1a10.ram_block_type = "auto";

cyclonev_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(rden_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a6.clk0_core_clock_enable = "ena0";
defparam ram_block1a6.clk1_core_clock_enable = "ena1";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "processor_cpu:cpu|processor_cpu_ic_data_module:processor_cpu_ic_data|altsyncram:the_altsyncram|altsyncram_ekj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 9;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 511;
defparam ram_block1a6.port_a_logical_ram_depth = 512;
defparam ram_block1a6.port_a_logical_ram_width = 32;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_address_clear = "none";
defparam ram_block1a6.port_b_address_clock = "clock1";
defparam ram_block1a6.port_b_address_width = 9;
defparam ram_block1a6.port_b_data_out_clear = "none";
defparam ram_block1a6.port_b_data_out_clock = "none";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 511;
defparam ram_block1a6.port_b_logical_ram_depth = 512;
defparam ram_block1a6.port_b_logical_ram_width = 32;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock1";
defparam ram_block1a6.ram_block_type = "auto";

cyclonev_ram_block ram_block1a8(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(rden_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a8_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a8.clk0_core_clock_enable = "ena0";
defparam ram_block1a8.clk1_core_clock_enable = "ena1";
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.logical_ram_name = "processor_cpu:cpu|processor_cpu_ic_data_module:processor_cpu_ic_data|altsyncram:the_altsyncram|altsyncram_ekj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a8.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a8.operation_mode = "dual_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 9;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 511;
defparam ram_block1a8.port_a_logical_ram_depth = 512;
defparam ram_block1a8.port_a_logical_ram_width = 32;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a8.port_b_address_clear = "none";
defparam ram_block1a8.port_b_address_clock = "clock1";
defparam ram_block1a8.port_b_address_width = 9;
defparam ram_block1a8.port_b_data_out_clear = "none";
defparam ram_block1a8.port_b_data_out_clock = "none";
defparam ram_block1a8.port_b_data_width = 1;
defparam ram_block1a8.port_b_first_address = 0;
defparam ram_block1a8.port_b_first_bit_number = 8;
defparam ram_block1a8.port_b_last_address = 511;
defparam ram_block1a8.port_b_logical_ram_depth = 512;
defparam ram_block1a8.port_b_logical_ram_width = 32;
defparam ram_block1a8.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a8.port_b_read_enable_clock = "clock1";
defparam ram_block1a8.ram_block_type = "auto";

cyclonev_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(rden_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a7.clk0_core_clock_enable = "ena0";
defparam ram_block1a7.clk1_core_clock_enable = "ena1";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "processor_cpu:cpu|processor_cpu_ic_data_module:processor_cpu_ic_data|altsyncram:the_altsyncram|altsyncram_ekj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 9;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 511;
defparam ram_block1a7.port_a_logical_ram_depth = 512;
defparam ram_block1a7.port_a_logical_ram_width = 32;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_address_clear = "none";
defparam ram_block1a7.port_b_address_clock = "clock1";
defparam ram_block1a7.port_b_address_width = 9;
defparam ram_block1a7.port_b_data_out_clear = "none";
defparam ram_block1a7.port_b_data_out_clock = "none";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 511;
defparam ram_block1a7.port_b_logical_ram_depth = 512;
defparam ram_block1a7.port_b_logical_ram_width = 32;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock1";
defparam ram_block1a7.ram_block_type = "auto";

cyclonev_ram_block ram_block1a20(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(rden_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[20]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a20_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a20.clk0_core_clock_enable = "ena0";
defparam ram_block1a20.clk1_core_clock_enable = "ena1";
defparam ram_block1a20.data_interleave_offset_in_bits = 1;
defparam ram_block1a20.data_interleave_width_in_bits = 1;
defparam ram_block1a20.logical_ram_name = "processor_cpu:cpu|processor_cpu_ic_data_module:processor_cpu_ic_data|altsyncram:the_altsyncram|altsyncram_ekj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a20.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a20.operation_mode = "dual_port";
defparam ram_block1a20.port_a_address_clear = "none";
defparam ram_block1a20.port_a_address_width = 9;
defparam ram_block1a20.port_a_data_out_clear = "none";
defparam ram_block1a20.port_a_data_out_clock = "none";
defparam ram_block1a20.port_a_data_width = 1;
defparam ram_block1a20.port_a_first_address = 0;
defparam ram_block1a20.port_a_first_bit_number = 20;
defparam ram_block1a20.port_a_last_address = 511;
defparam ram_block1a20.port_a_logical_ram_depth = 512;
defparam ram_block1a20.port_a_logical_ram_width = 32;
defparam ram_block1a20.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a20.port_b_address_clear = "none";
defparam ram_block1a20.port_b_address_clock = "clock1";
defparam ram_block1a20.port_b_address_width = 9;
defparam ram_block1a20.port_b_data_out_clear = "none";
defparam ram_block1a20.port_b_data_out_clock = "none";
defparam ram_block1a20.port_b_data_width = 1;
defparam ram_block1a20.port_b_first_address = 0;
defparam ram_block1a20.port_b_first_bit_number = 20;
defparam ram_block1a20.port_b_last_address = 511;
defparam ram_block1a20.port_b_logical_ram_depth = 512;
defparam ram_block1a20.port_b_logical_ram_width = 32;
defparam ram_block1a20.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a20.port_b_read_enable_clock = "clock1";
defparam ram_block1a20.ram_block_type = "auto";

cyclonev_ram_block ram_block1a19(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(rden_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[19]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a19_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a19.clk0_core_clock_enable = "ena0";
defparam ram_block1a19.clk1_core_clock_enable = "ena1";
defparam ram_block1a19.data_interleave_offset_in_bits = 1;
defparam ram_block1a19.data_interleave_width_in_bits = 1;
defparam ram_block1a19.logical_ram_name = "processor_cpu:cpu|processor_cpu_ic_data_module:processor_cpu_ic_data|altsyncram:the_altsyncram|altsyncram_ekj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a19.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a19.operation_mode = "dual_port";
defparam ram_block1a19.port_a_address_clear = "none";
defparam ram_block1a19.port_a_address_width = 9;
defparam ram_block1a19.port_a_data_out_clear = "none";
defparam ram_block1a19.port_a_data_out_clock = "none";
defparam ram_block1a19.port_a_data_width = 1;
defparam ram_block1a19.port_a_first_address = 0;
defparam ram_block1a19.port_a_first_bit_number = 19;
defparam ram_block1a19.port_a_last_address = 511;
defparam ram_block1a19.port_a_logical_ram_depth = 512;
defparam ram_block1a19.port_a_logical_ram_width = 32;
defparam ram_block1a19.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a19.port_b_address_clear = "none";
defparam ram_block1a19.port_b_address_clock = "clock1";
defparam ram_block1a19.port_b_address_width = 9;
defparam ram_block1a19.port_b_data_out_clear = "none";
defparam ram_block1a19.port_b_data_out_clock = "none";
defparam ram_block1a19.port_b_data_width = 1;
defparam ram_block1a19.port_b_first_address = 0;
defparam ram_block1a19.port_b_first_bit_number = 19;
defparam ram_block1a19.port_b_last_address = 511;
defparam ram_block1a19.port_b_logical_ram_depth = 512;
defparam ram_block1a19.port_b_logical_ram_width = 32;
defparam ram_block1a19.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a19.port_b_read_enable_clock = "clock1";
defparam ram_block1a19.ram_block_type = "auto";

cyclonev_ram_block ram_block1a18(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(rden_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[18]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a18_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a18.clk0_core_clock_enable = "ena0";
defparam ram_block1a18.clk1_core_clock_enable = "ena1";
defparam ram_block1a18.data_interleave_offset_in_bits = 1;
defparam ram_block1a18.data_interleave_width_in_bits = 1;
defparam ram_block1a18.logical_ram_name = "processor_cpu:cpu|processor_cpu_ic_data_module:processor_cpu_ic_data|altsyncram:the_altsyncram|altsyncram_ekj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a18.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a18.operation_mode = "dual_port";
defparam ram_block1a18.port_a_address_clear = "none";
defparam ram_block1a18.port_a_address_width = 9;
defparam ram_block1a18.port_a_data_out_clear = "none";
defparam ram_block1a18.port_a_data_out_clock = "none";
defparam ram_block1a18.port_a_data_width = 1;
defparam ram_block1a18.port_a_first_address = 0;
defparam ram_block1a18.port_a_first_bit_number = 18;
defparam ram_block1a18.port_a_last_address = 511;
defparam ram_block1a18.port_a_logical_ram_depth = 512;
defparam ram_block1a18.port_a_logical_ram_width = 32;
defparam ram_block1a18.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a18.port_b_address_clear = "none";
defparam ram_block1a18.port_b_address_clock = "clock1";
defparam ram_block1a18.port_b_address_width = 9;
defparam ram_block1a18.port_b_data_out_clear = "none";
defparam ram_block1a18.port_b_data_out_clock = "none";
defparam ram_block1a18.port_b_data_width = 1;
defparam ram_block1a18.port_b_first_address = 0;
defparam ram_block1a18.port_b_first_bit_number = 18;
defparam ram_block1a18.port_b_last_address = 511;
defparam ram_block1a18.port_b_logical_ram_depth = 512;
defparam ram_block1a18.port_b_logical_ram_width = 32;
defparam ram_block1a18.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a18.port_b_read_enable_clock = "clock1";
defparam ram_block1a18.ram_block_type = "auto";

cyclonev_ram_block ram_block1a17(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(rden_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[17]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a17_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a17.clk0_core_clock_enable = "ena0";
defparam ram_block1a17.clk1_core_clock_enable = "ena1";
defparam ram_block1a17.data_interleave_offset_in_bits = 1;
defparam ram_block1a17.data_interleave_width_in_bits = 1;
defparam ram_block1a17.logical_ram_name = "processor_cpu:cpu|processor_cpu_ic_data_module:processor_cpu_ic_data|altsyncram:the_altsyncram|altsyncram_ekj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a17.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a17.operation_mode = "dual_port";
defparam ram_block1a17.port_a_address_clear = "none";
defparam ram_block1a17.port_a_address_width = 9;
defparam ram_block1a17.port_a_data_out_clear = "none";
defparam ram_block1a17.port_a_data_out_clock = "none";
defparam ram_block1a17.port_a_data_width = 1;
defparam ram_block1a17.port_a_first_address = 0;
defparam ram_block1a17.port_a_first_bit_number = 17;
defparam ram_block1a17.port_a_last_address = 511;
defparam ram_block1a17.port_a_logical_ram_depth = 512;
defparam ram_block1a17.port_a_logical_ram_width = 32;
defparam ram_block1a17.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a17.port_b_address_clear = "none";
defparam ram_block1a17.port_b_address_clock = "clock1";
defparam ram_block1a17.port_b_address_width = 9;
defparam ram_block1a17.port_b_data_out_clear = "none";
defparam ram_block1a17.port_b_data_out_clock = "none";
defparam ram_block1a17.port_b_data_width = 1;
defparam ram_block1a17.port_b_first_address = 0;
defparam ram_block1a17.port_b_first_bit_number = 17;
defparam ram_block1a17.port_b_last_address = 511;
defparam ram_block1a17.port_b_logical_ram_depth = 512;
defparam ram_block1a17.port_b_logical_ram_width = 32;
defparam ram_block1a17.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a17.port_b_read_enable_clock = "clock1";
defparam ram_block1a17.ram_block_type = "auto";

cyclonev_ram_block ram_block1a9(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(rden_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a9_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a9.clk0_core_clock_enable = "ena0";
defparam ram_block1a9.clk1_core_clock_enable = "ena1";
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.logical_ram_name = "processor_cpu:cpu|processor_cpu_ic_data_module:processor_cpu_ic_data|altsyncram:the_altsyncram|altsyncram_ekj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a9.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a9.operation_mode = "dual_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 9;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 511;
defparam ram_block1a9.port_a_logical_ram_depth = 512;
defparam ram_block1a9.port_a_logical_ram_width = 32;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a9.port_b_address_clear = "none";
defparam ram_block1a9.port_b_address_clock = "clock1";
defparam ram_block1a9.port_b_address_width = 9;
defparam ram_block1a9.port_b_data_out_clear = "none";
defparam ram_block1a9.port_b_data_out_clock = "none";
defparam ram_block1a9.port_b_data_width = 1;
defparam ram_block1a9.port_b_first_address = 0;
defparam ram_block1a9.port_b_first_bit_number = 9;
defparam ram_block1a9.port_b_last_address = 511;
defparam ram_block1a9.port_b_logical_ram_depth = 512;
defparam ram_block1a9.port_b_logical_ram_width = 32;
defparam ram_block1a9.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a9.port_b_read_enable_clock = "clock1";
defparam ram_block1a9.ram_block_type = "auto";

endmodule

module processor_processor_cpu_ic_tag_module (
	q_b_5,
	q_b_1,
	q_b_4,
	q_b_0,
	q_b_2,
	q_b_3,
	q_b_11,
	q_b_13,
	q_b_10,
	q_b_12,
	ic_tag_wraddress_0,
	ic_fill_valid_bits_5,
	ic_fill_valid_bits_7,
	ic_fill_valid_bits_4,
	q_b_7,
	q_b_9,
	q_b_6,
	q_b_8,
	ic_fill_valid_bits_6,
	ic_fill_valid_bits_1,
	ic_fill_valid_bits_3,
	ic_fill_valid_bits_0,
	ic_fill_valid_bits_2,
	W_stall,
	ic_fill_tag_5,
	ic_fill_tag_4,
	ic_fill_tag_3,
	ic_fill_tag_2,
	ic_fill_tag_1,
	ic_fill_tag_0,
	F_ic_tag_rd_addr_nxt_0,
	F_ic_tag_rd_addr_nxt_1,
	F_ic_tag_rd_addr_nxt_2,
	F_ic_tag_rd_addr_nxt_3,
	F_ic_tag_rd_addr_nxt_4,
	F_ic_tag_rd_addr_nxt_5,
	ic_tag_wren,
	ic_tag_wraddress_1,
	ic_tag_wraddress_2,
	ic_tag_wraddress_3,
	ic_tag_wraddress_4,
	ic_tag_wraddress_5,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_5;
output 	q_b_1;
output 	q_b_4;
output 	q_b_0;
output 	q_b_2;
output 	q_b_3;
output 	q_b_11;
output 	q_b_13;
output 	q_b_10;
output 	q_b_12;
input 	ic_tag_wraddress_0;
input 	ic_fill_valid_bits_5;
input 	ic_fill_valid_bits_7;
input 	ic_fill_valid_bits_4;
output 	q_b_7;
output 	q_b_9;
output 	q_b_6;
output 	q_b_8;
input 	ic_fill_valid_bits_6;
input 	ic_fill_valid_bits_1;
input 	ic_fill_valid_bits_3;
input 	ic_fill_valid_bits_0;
input 	ic_fill_valid_bits_2;
input 	W_stall;
input 	ic_fill_tag_5;
input 	ic_fill_tag_4;
input 	ic_fill_tag_3;
input 	ic_fill_tag_2;
input 	ic_fill_tag_1;
input 	ic_fill_tag_0;
input 	F_ic_tag_rd_addr_nxt_0;
input 	F_ic_tag_rd_addr_nxt_1;
input 	F_ic_tag_rd_addr_nxt_2;
input 	F_ic_tag_rd_addr_nxt_3;
input 	F_ic_tag_rd_addr_nxt_4;
input 	F_ic_tag_rd_addr_nxt_5;
input 	ic_tag_wren;
input 	ic_tag_wraddress_1;
input 	ic_tag_wraddress_2;
input 	ic_tag_wraddress_3;
input 	ic_tag_wraddress_4;
input 	ic_tag_wraddress_5;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



processor_altsyncram_2 the_altsyncram(
	.q_b({q_b_unconnected_wire_31,q_b_unconnected_wire_30,q_b_unconnected_wire_29,q_b_unconnected_wire_28,q_b_unconnected_wire_27,q_b_unconnected_wire_26,q_b_unconnected_wire_25,q_b_unconnected_wire_24,q_b_unconnected_wire_23,q_b_unconnected_wire_22,q_b_unconnected_wire_21,
q_b_unconnected_wire_20,q_b_unconnected_wire_19,q_b_unconnected_wire_18,q_b_unconnected_wire_17,q_b_unconnected_wire_16,q_b_unconnected_wire_15,q_b_unconnected_wire_14,q_b_13,q_b_12,q_b_11,q_b_10,q_b_9,q_b_8,q_b_7,q_b_6,q_b_5,q_b_4,q_b_3,q_b_2,q_b_1,q_b_0}),
	.address_a({gnd,gnd,gnd,gnd,gnd,gnd,gnd,ic_tag_wraddress_5,ic_tag_wraddress_4,ic_tag_wraddress_3,ic_tag_wraddress_2,ic_tag_wraddress_1,ic_tag_wraddress_0}),
	.data_a({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,ic_fill_valid_bits_7,ic_fill_valid_bits_6,ic_fill_valid_bits_5,ic_fill_valid_bits_4,ic_fill_valid_bits_3,ic_fill_valid_bits_2,ic_fill_valid_bits_1,ic_fill_valid_bits_0,ic_fill_tag_5,ic_fill_tag_4,ic_fill_tag_3,
ic_fill_tag_2,ic_fill_tag_1,ic_fill_tag_0}),
	.rden_b(W_stall),
	.address_b({gnd,gnd,gnd,F_ic_tag_rd_addr_nxt_5,F_ic_tag_rd_addr_nxt_4,F_ic_tag_rd_addr_nxt_3,F_ic_tag_rd_addr_nxt_2,F_ic_tag_rd_addr_nxt_1,F_ic_tag_rd_addr_nxt_0}),
	.wren_a(ic_tag_wren),
	.clock0(clk_clk));

endmodule

module processor_altsyncram_2 (
	q_b,
	address_a,
	data_a,
	rden_b,
	address_b,
	wren_a,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[31:0] q_b;
input 	[12:0] address_a;
input 	[31:0] data_a;
input 	rden_b;
input 	[8:0] address_b;
input 	wren_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



processor_altsyncram_van1 auto_generated(
	.q_b({q_b[13],q_b[12],q_b[11],q_b[10],q_b[9],q_b[8],q_b[7],q_b[6],q_b[5],q_b[4],q_b[3],q_b[2],q_b[1],q_b[0]}),
	.address_a({address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.data_a({data_a[13],data_a[12],data_a[11],data_a[10],data_a[9],data_a[8],data_a[7],data_a[6],data_a[5],data_a[4],data_a[3],data_a[2],data_a[1],data_a[0]}),
	.rden_b(rden_b),
	.address_b({address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.wren_a(wren_a),
	.clock0(clock0));

endmodule

module processor_altsyncram_van1 (
	q_b,
	address_a,
	data_a,
	rden_b,
	address_b,
	wren_a,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[13:0] q_b;
input 	[5:0] address_a;
input 	[13:0] data_a;
input 	rden_b;
input 	[5:0] address_b;
input 	wren_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a1_PORTBDATAOUT_bus;
wire [143:0] ram_block1a4_PORTBDATAOUT_bus;
wire [143:0] ram_block1a0_PORTBDATAOUT_bus;
wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;
wire [143:0] ram_block1a11_PORTBDATAOUT_bus;
wire [143:0] ram_block1a13_PORTBDATAOUT_bus;
wire [143:0] ram_block1a10_PORTBDATAOUT_bus;
wire [143:0] ram_block1a12_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a9_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a8_PORTBDATAOUT_bus;

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

assign q_b[2] = ram_block1a2_PORTBDATAOUT_bus[0];

assign q_b[3] = ram_block1a3_PORTBDATAOUT_bus[0];

assign q_b[11] = ram_block1a11_PORTBDATAOUT_bus[0];

assign q_b[13] = ram_block1a13_PORTBDATAOUT_bus[0];

assign q_b[10] = ram_block1a10_PORTBDATAOUT_bus[0];

assign q_b[12] = ram_block1a12_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_b[9] = ram_block1a9_PORTBDATAOUT_bus[0];

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_b[8] = ram_block1a8_PORTBDATAOUT_bus[0];

cyclonev_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.init_file = "processor_cpu_ic_tag_ram.mif";
defparam ram_block1a5.init_file_layout = "port_b";
defparam ram_block1a5.logical_ram_name = "processor_cpu:cpu|processor_cpu_ic_tag_module:processor_cpu_ic_tag|altsyncram:the_altsyncram|altsyncram_van1:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "old";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 6;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 63;
defparam ram_block1a5.port_a_logical_ram_depth = 64;
defparam ram_block1a5.port_a_logical_ram_width = 14;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_address_clear = "none";
defparam ram_block1a5.port_b_address_clock = "clock0";
defparam ram_block1a5.port_b_address_width = 6;
defparam ram_block1a5.port_b_data_out_clear = "none";
defparam ram_block1a5.port_b_data_out_clock = "none";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 63;
defparam ram_block1a5.port_b_logical_ram_depth = 64;
defparam ram_block1a5.port_b_logical_ram_width = 14;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock0";
defparam ram_block1a5.ram_block_type = "auto";
defparam ram_block1a5.mem_init0 = "7209A6A81568A156";

cyclonev_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.init_file = "processor_cpu_ic_tag_ram.mif";
defparam ram_block1a1.init_file_layout = "port_b";
defparam ram_block1a1.logical_ram_name = "processor_cpu:cpu|processor_cpu_ic_tag_module:processor_cpu_ic_tag|altsyncram:the_altsyncram|altsyncram_van1:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "old";
defparam ram_block1a1.operation_mode = "dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 6;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 63;
defparam ram_block1a1.port_a_logical_ram_depth = 64;
defparam ram_block1a1.port_a_logical_ram_width = 14;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_address_clear = "none";
defparam ram_block1a1.port_b_address_clock = "clock0";
defparam ram_block1a1.port_b_address_width = 6;
defparam ram_block1a1.port_b_data_out_clear = "none";
defparam ram_block1a1.port_b_data_out_clock = "none";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 63;
defparam ram_block1a1.port_b_logical_ram_depth = 64;
defparam ram_block1a1.port_b_logical_ram_width = 14;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock0";
defparam ram_block1a1.ram_block_type = "auto";
defparam ram_block1a1.mem_init0 = "198D03846DA98D04";

cyclonev_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.init_file = "processor_cpu_ic_tag_ram.mif";
defparam ram_block1a4.init_file_layout = "port_b";
defparam ram_block1a4.logical_ram_name = "processor_cpu:cpu|processor_cpu_ic_tag_module:processor_cpu_ic_tag|altsyncram:the_altsyncram|altsyncram_van1:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "old";
defparam ram_block1a4.operation_mode = "dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 6;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 63;
defparam ram_block1a4.port_a_logical_ram_depth = 64;
defparam ram_block1a4.port_a_logical_ram_width = 14;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_address_clear = "none";
defparam ram_block1a4.port_b_address_clock = "clock0";
defparam ram_block1a4.port_b_address_width = 6;
defparam ram_block1a4.port_b_data_out_clear = "none";
defparam ram_block1a4.port_b_data_out_clock = "none";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 63;
defparam ram_block1a4.port_b_logical_ram_depth = 64;
defparam ram_block1a4.port_b_logical_ram_width = 14;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock0";
defparam ram_block1a4.ram_block_type = "auto";
defparam ram_block1a4.mem_init0 = "C7150B3DCE44583B";

cyclonev_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.init_file = "processor_cpu_ic_tag_ram.mif";
defparam ram_block1a0.init_file_layout = "port_b";
defparam ram_block1a0.logical_ram_name = "processor_cpu:cpu|processor_cpu_ic_tag_module:processor_cpu_ic_tag|altsyncram:the_altsyncram|altsyncram_van1:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "old";
defparam ram_block1a0.operation_mode = "dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 6;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 63;
defparam ram_block1a0.port_a_logical_ram_depth = 64;
defparam ram_block1a0.port_a_logical_ram_width = 14;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_address_clear = "none";
defparam ram_block1a0.port_b_address_clock = "clock0";
defparam ram_block1a0.port_b_address_width = 6;
defparam ram_block1a0.port_b_data_out_clear = "none";
defparam ram_block1a0.port_b_data_out_clock = "none";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 63;
defparam ram_block1a0.port_b_logical_ram_depth = 64;
defparam ram_block1a0.port_b_logical_ram_width = 14;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock0";
defparam ram_block1a0.ram_block_type = "auto";
defparam ram_block1a0.mem_init0 = "B4E2FBAE751F1E7B";

cyclonev_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.init_file = "processor_cpu_ic_tag_ram.mif";
defparam ram_block1a2.init_file_layout = "port_b";
defparam ram_block1a2.logical_ram_name = "processor_cpu:cpu|processor_cpu_ic_tag_module:processor_cpu_ic_tag|altsyncram:the_altsyncram|altsyncram_van1:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "old";
defparam ram_block1a2.operation_mode = "dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 6;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 63;
defparam ram_block1a2.port_a_logical_ram_depth = 64;
defparam ram_block1a2.port_a_logical_ram_width = 14;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_address_clear = "none";
defparam ram_block1a2.port_b_address_clock = "clock0";
defparam ram_block1a2.port_b_address_width = 6;
defparam ram_block1a2.port_b_data_out_clear = "none";
defparam ram_block1a2.port_b_data_out_clock = "none";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 63;
defparam ram_block1a2.port_b_logical_ram_depth = 64;
defparam ram_block1a2.port_b_logical_ram_width = 14;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock0";
defparam ram_block1a2.ram_block_type = "auto";
defparam ram_block1a2.mem_init0 = "66F33435CC960198";

cyclonev_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.init_file = "processor_cpu_ic_tag_ram.mif";
defparam ram_block1a3.init_file_layout = "port_b";
defparam ram_block1a3.logical_ram_name = "processor_cpu:cpu|processor_cpu_ic_tag_module:processor_cpu_ic_tag|altsyncram:the_altsyncram|altsyncram_van1:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "old";
defparam ram_block1a3.operation_mode = "dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 6;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 63;
defparam ram_block1a3.port_a_logical_ram_depth = 64;
defparam ram_block1a3.port_a_logical_ram_width = 14;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_address_clear = "none";
defparam ram_block1a3.port_b_address_clock = "clock0";
defparam ram_block1a3.port_b_address_width = 6;
defparam ram_block1a3.port_b_data_out_clear = "none";
defparam ram_block1a3.port_b_data_out_clock = "none";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 63;
defparam ram_block1a3.port_b_logical_ram_depth = 64;
defparam ram_block1a3.port_b_logical_ram_width = 14;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock0";
defparam ram_block1a3.ram_block_type = "auto";
defparam ram_block1a3.mem_init0 = "32C19C540815BA17";

cyclonev_ram_block ram_block1a11(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a11_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.init_file = "processor_cpu_ic_tag_ram.mif";
defparam ram_block1a11.init_file_layout = "port_b";
defparam ram_block1a11.logical_ram_name = "processor_cpu:cpu|processor_cpu_ic_tag_module:processor_cpu_ic_tag|altsyncram:the_altsyncram|altsyncram_van1:auto_generated|ALTSYNCRAM";
defparam ram_block1a11.mixed_port_feed_through_mode = "old";
defparam ram_block1a11.operation_mode = "dual_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 6;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 63;
defparam ram_block1a11.port_a_logical_ram_depth = 64;
defparam ram_block1a11.port_a_logical_ram_width = 14;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a11.port_b_address_clear = "none";
defparam ram_block1a11.port_b_address_clock = "clock0";
defparam ram_block1a11.port_b_address_width = 6;
defparam ram_block1a11.port_b_data_out_clear = "none";
defparam ram_block1a11.port_b_data_out_clock = "none";
defparam ram_block1a11.port_b_data_width = 1;
defparam ram_block1a11.port_b_first_address = 0;
defparam ram_block1a11.port_b_first_bit_number = 11;
defparam ram_block1a11.port_b_last_address = 63;
defparam ram_block1a11.port_b_logical_ram_depth = 64;
defparam ram_block1a11.port_b_logical_ram_width = 14;
defparam ram_block1a11.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a11.port_b_read_enable_clock = "clock0";
defparam ram_block1a11.ram_block_type = "auto";
defparam ram_block1a11.mem_init0 = "864713E5C66BCE07";

cyclonev_ram_block ram_block1a13(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a13_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.init_file = "processor_cpu_ic_tag_ram.mif";
defparam ram_block1a13.init_file_layout = "port_b";
defparam ram_block1a13.logical_ram_name = "processor_cpu:cpu|processor_cpu_ic_tag_module:processor_cpu_ic_tag|altsyncram:the_altsyncram|altsyncram_van1:auto_generated|ALTSYNCRAM";
defparam ram_block1a13.mixed_port_feed_through_mode = "old";
defparam ram_block1a13.operation_mode = "dual_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 6;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 63;
defparam ram_block1a13.port_a_logical_ram_depth = 64;
defparam ram_block1a13.port_a_logical_ram_width = 14;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a13.port_b_address_clear = "none";
defparam ram_block1a13.port_b_address_clock = "clock0";
defparam ram_block1a13.port_b_address_width = 6;
defparam ram_block1a13.port_b_data_out_clear = "none";
defparam ram_block1a13.port_b_data_out_clock = "none";
defparam ram_block1a13.port_b_data_width = 1;
defparam ram_block1a13.port_b_first_address = 0;
defparam ram_block1a13.port_b_first_bit_number = 13;
defparam ram_block1a13.port_b_last_address = 63;
defparam ram_block1a13.port_b_logical_ram_depth = 64;
defparam ram_block1a13.port_b_logical_ram_width = 14;
defparam ram_block1a13.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a13.port_b_read_enable_clock = "clock0";
defparam ram_block1a13.ram_block_type = "auto";
defparam ram_block1a13.mem_init0 = "E0EC38012A3EDBCD";

cyclonev_ram_block ram_block1a10(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a10_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.init_file = "processor_cpu_ic_tag_ram.mif";
defparam ram_block1a10.init_file_layout = "port_b";
defparam ram_block1a10.logical_ram_name = "processor_cpu:cpu|processor_cpu_ic_tag_module:processor_cpu_ic_tag|altsyncram:the_altsyncram|altsyncram_van1:auto_generated|ALTSYNCRAM";
defparam ram_block1a10.mixed_port_feed_through_mode = "old";
defparam ram_block1a10.operation_mode = "dual_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 6;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 63;
defparam ram_block1a10.port_a_logical_ram_depth = 64;
defparam ram_block1a10.port_a_logical_ram_width = 14;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a10.port_b_address_clear = "none";
defparam ram_block1a10.port_b_address_clock = "clock0";
defparam ram_block1a10.port_b_address_width = 6;
defparam ram_block1a10.port_b_data_out_clear = "none";
defparam ram_block1a10.port_b_data_out_clock = "none";
defparam ram_block1a10.port_b_data_width = 1;
defparam ram_block1a10.port_b_first_address = 0;
defparam ram_block1a10.port_b_first_bit_number = 10;
defparam ram_block1a10.port_b_last_address = 63;
defparam ram_block1a10.port_b_logical_ram_depth = 64;
defparam ram_block1a10.port_b_logical_ram_width = 14;
defparam ram_block1a10.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a10.port_b_read_enable_clock = "clock0";
defparam ram_block1a10.ram_block_type = "auto";
defparam ram_block1a10.mem_init0 = "B7985C4CB0BBC968";

cyclonev_ram_block ram_block1a12(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a12_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.init_file = "processor_cpu_ic_tag_ram.mif";
defparam ram_block1a12.init_file_layout = "port_b";
defparam ram_block1a12.logical_ram_name = "processor_cpu:cpu|processor_cpu_ic_tag_module:processor_cpu_ic_tag|altsyncram:the_altsyncram|altsyncram_van1:auto_generated|ALTSYNCRAM";
defparam ram_block1a12.mixed_port_feed_through_mode = "old";
defparam ram_block1a12.operation_mode = "dual_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 6;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 63;
defparam ram_block1a12.port_a_logical_ram_depth = 64;
defparam ram_block1a12.port_a_logical_ram_width = 14;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a12.port_b_address_clear = "none";
defparam ram_block1a12.port_b_address_clock = "clock0";
defparam ram_block1a12.port_b_address_width = 6;
defparam ram_block1a12.port_b_data_out_clear = "none";
defparam ram_block1a12.port_b_data_out_clock = "none";
defparam ram_block1a12.port_b_data_width = 1;
defparam ram_block1a12.port_b_first_address = 0;
defparam ram_block1a12.port_b_first_bit_number = 12;
defparam ram_block1a12.port_b_last_address = 63;
defparam ram_block1a12.port_b_logical_ram_depth = 64;
defparam ram_block1a12.port_b_logical_ram_width = 14;
defparam ram_block1a12.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a12.port_b_read_enable_clock = "clock0";
defparam ram_block1a12.ram_block_type = "auto";
defparam ram_block1a12.mem_init0 = "F35ABCDC9F60190A";

cyclonev_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.init_file = "processor_cpu_ic_tag_ram.mif";
defparam ram_block1a7.init_file_layout = "port_b";
defparam ram_block1a7.logical_ram_name = "processor_cpu:cpu|processor_cpu_ic_tag_module:processor_cpu_ic_tag|altsyncram:the_altsyncram|altsyncram_van1:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "old";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 6;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 63;
defparam ram_block1a7.port_a_logical_ram_depth = 64;
defparam ram_block1a7.port_a_logical_ram_width = 14;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_address_clear = "none";
defparam ram_block1a7.port_b_address_clock = "clock0";
defparam ram_block1a7.port_b_address_width = 6;
defparam ram_block1a7.port_b_data_out_clear = "none";
defparam ram_block1a7.port_b_data_out_clock = "none";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 63;
defparam ram_block1a7.port_b_logical_ram_depth = 64;
defparam ram_block1a7.port_b_logical_ram_width = 14;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock0";
defparam ram_block1a7.ram_block_type = "auto";
defparam ram_block1a7.mem_init0 = "40349E904F8351BF";

cyclonev_ram_block ram_block1a9(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a9_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.init_file = "processor_cpu_ic_tag_ram.mif";
defparam ram_block1a9.init_file_layout = "port_b";
defparam ram_block1a9.logical_ram_name = "processor_cpu:cpu|processor_cpu_ic_tag_module:processor_cpu_ic_tag|altsyncram:the_altsyncram|altsyncram_van1:auto_generated|ALTSYNCRAM";
defparam ram_block1a9.mixed_port_feed_through_mode = "old";
defparam ram_block1a9.operation_mode = "dual_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 6;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 63;
defparam ram_block1a9.port_a_logical_ram_depth = 64;
defparam ram_block1a9.port_a_logical_ram_width = 14;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a9.port_b_address_clear = "none";
defparam ram_block1a9.port_b_address_clock = "clock0";
defparam ram_block1a9.port_b_address_width = 6;
defparam ram_block1a9.port_b_data_out_clear = "none";
defparam ram_block1a9.port_b_data_out_clock = "none";
defparam ram_block1a9.port_b_data_width = 1;
defparam ram_block1a9.port_b_first_address = 0;
defparam ram_block1a9.port_b_first_bit_number = 9;
defparam ram_block1a9.port_b_last_address = 63;
defparam ram_block1a9.port_b_logical_ram_depth = 64;
defparam ram_block1a9.port_b_logical_ram_width = 14;
defparam ram_block1a9.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a9.port_b_read_enable_clock = "clock0";
defparam ram_block1a9.ram_block_type = "auto";
defparam ram_block1a9.mem_init0 = "0D6F81A0DC328FD6";

cyclonev_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.init_file = "processor_cpu_ic_tag_ram.mif";
defparam ram_block1a6.init_file_layout = "port_b";
defparam ram_block1a6.logical_ram_name = "processor_cpu:cpu|processor_cpu_ic_tag_module:processor_cpu_ic_tag|altsyncram:the_altsyncram|altsyncram_van1:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "old";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 6;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 63;
defparam ram_block1a6.port_a_logical_ram_depth = 64;
defparam ram_block1a6.port_a_logical_ram_width = 14;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_address_clear = "none";
defparam ram_block1a6.port_b_address_clock = "clock0";
defparam ram_block1a6.port_b_address_width = 6;
defparam ram_block1a6.port_b_data_out_clear = "none";
defparam ram_block1a6.port_b_data_out_clock = "none";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 63;
defparam ram_block1a6.port_b_logical_ram_depth = 64;
defparam ram_block1a6.port_b_logical_ram_width = 14;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock0";
defparam ram_block1a6.ram_block_type = "auto";
defparam ram_block1a6.mem_init0 = "4F2996DA16385CF2";

cyclonev_ram_block ram_block1a8(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a8_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.init_file = "processor_cpu_ic_tag_ram.mif";
defparam ram_block1a8.init_file_layout = "port_b";
defparam ram_block1a8.logical_ram_name = "processor_cpu:cpu|processor_cpu_ic_tag_module:processor_cpu_ic_tag|altsyncram:the_altsyncram|altsyncram_van1:auto_generated|ALTSYNCRAM";
defparam ram_block1a8.mixed_port_feed_through_mode = "old";
defparam ram_block1a8.operation_mode = "dual_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 6;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 63;
defparam ram_block1a8.port_a_logical_ram_depth = 64;
defparam ram_block1a8.port_a_logical_ram_width = 14;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a8.port_b_address_clear = "none";
defparam ram_block1a8.port_b_address_clock = "clock0";
defparam ram_block1a8.port_b_address_width = 6;
defparam ram_block1a8.port_b_data_out_clear = "none";
defparam ram_block1a8.port_b_data_out_clock = "none";
defparam ram_block1a8.port_b_data_width = 1;
defparam ram_block1a8.port_b_first_address = 0;
defparam ram_block1a8.port_b_first_bit_number = 8;
defparam ram_block1a8.port_b_last_address = 63;
defparam ram_block1a8.port_b_logical_ram_depth = 64;
defparam ram_block1a8.port_b_logical_ram_width = 14;
defparam ram_block1a8.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a8.port_b_read_enable_clock = "clock0";
defparam ram_block1a8.ram_block_type = "auto";
defparam ram_block1a8.mem_init0 = "F63F2250392C148C";

endmodule

module processor_processor_cpu_nios2_oci (
	readdata_0,
	readdata_16,
	readdata_8,
	readdata_24,
	readdata_5,
	readdata_21,
	readdata_13,
	readdata_29,
	readdata_4,
	readdata_20,
	readdata_12,
	readdata_28,
	readdata_6,
	readdata_22,
	readdata_14,
	readdata_30,
	readdata_7,
	readdata_23,
	readdata_15,
	readdata_31,
	readdata_11,
	readdata_27,
	readdata_10,
	readdata_26,
	readdata_25,
	readdata_9,
	readdata_3,
	readdata_19,
	readdata_2,
	readdata_18,
	readdata_1,
	readdata_17,
	sr_0,
	ir_out_0,
	ir_out_1,
	r_sync_rst,
	d_write,
	saved_grant_0,
	waitrequest,
	mem_used_1,
	hbreak_enabled,
	jtag_break,
	src2_valid,
	saved_grant_1,
	src0_valid,
	rf_source_valid,
	oci_single_step_mode,
	address_nxt,
	oci_ienable_16,
	r_early_rst,
	oci_ienable_1,
	writedata_nxt,
	debugaccess_nxt,
	byteenable_nxt,
	altera_internal_jtag,
	altera_internal_jtag1,
	state_1,
	state_4,
	virtual_ir_scan_reg,
	state_3,
	state_8,
	splitter_nodes_receive_1_3,
	irf_reg_0_2,
	irf_reg_1_2,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	readdata_0;
output 	readdata_16;
output 	readdata_8;
output 	readdata_24;
output 	readdata_5;
output 	readdata_21;
output 	readdata_13;
output 	readdata_29;
output 	readdata_4;
output 	readdata_20;
output 	readdata_12;
output 	readdata_28;
output 	readdata_6;
output 	readdata_22;
output 	readdata_14;
output 	readdata_30;
output 	readdata_7;
output 	readdata_23;
output 	readdata_15;
output 	readdata_31;
output 	readdata_11;
output 	readdata_27;
output 	readdata_10;
output 	readdata_26;
output 	readdata_25;
output 	readdata_9;
output 	readdata_3;
output 	readdata_19;
output 	readdata_2;
output 	readdata_18;
output 	readdata_1;
output 	readdata_17;
output 	sr_0;
output 	ir_out_0;
output 	ir_out_1;
input 	r_sync_rst;
input 	d_write;
input 	saved_grant_0;
output 	waitrequest;
input 	mem_used_1;
input 	hbreak_enabled;
output 	jtag_break;
input 	src2_valid;
input 	saved_grant_1;
input 	src0_valid;
input 	rf_source_valid;
output 	oci_single_step_mode;
input 	[8:0] address_nxt;
output 	oci_ienable_16;
input 	r_early_rst;
output 	oci_ienable_1;
input 	[31:0] writedata_nxt;
input 	debugaccess_nxt;
input 	[3:0] byteenable_nxt;
input 	altera_internal_jtag;
input 	altera_internal_jtag1;
input 	state_1;
input 	state_4;
input 	virtual_ir_scan_reg;
input 	state_3;
input 	state_8;
input 	splitter_nodes_receive_1_3;
input 	irf_reg_0_2;
input 	irf_reg_1_2;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \the_processor_cpu_nios2_oci_break|break_readreg[0]~q ;
wire \the_processor_cpu_nios2_oci_break|break_readreg[1]~q ;
wire \the_processor_cpu_nios2_ocimem|processor_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[0] ;
wire \the_processor_cpu_nios2_oci_break|break_readreg[2]~q ;
wire \the_processor_cpu_nios2_ocimem|MonDReg[2]~q ;
wire \the_processor_cpu_nios2_ocimem|processor_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[1] ;
wire \the_processor_cpu_nios2_oci_break|break_readreg[20]~q ;
wire \the_processor_cpu_nios2_ocimem|MonDReg[20]~q ;
wire \the_processor_cpu_nios2_oci_break|break_readreg[19]~q ;
wire \the_processor_cpu_nios2_ocimem|MonDReg[19]~q ;
wire \the_processor_cpu_nios2_oci_break|break_readreg[3]~q ;
wire \the_processor_cpu_nios2_ocimem|processor_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[2] ;
wire \the_processor_cpu_nios2_ocimem|processor_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[16] ;
wire \the_processor_cpu_nios2_ocimem|processor_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[8] ;
wire \the_processor_cpu_nios2_ocimem|processor_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[24] ;
wire \the_processor_cpu_nios2_oci_break|break_readreg[16]~q ;
wire \the_processor_cpu_nios2_ocimem|MonDReg[16]~q ;
wire \the_processor_cpu_nios2_oci_break|break_readreg[21]~q ;
wire \the_processor_cpu_nios2_ocimem|MonDReg[21]~q ;
wire \the_processor_cpu_nios2_ocimem|processor_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[20] ;
wire \the_processor_cpu_nios2_ocimem|processor_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[19] ;
wire \the_processor_cpu_nios2_oci_break|break_readreg[18]~q ;
wire \the_processor_cpu_nios2_oci_break|break_readreg[17]~q ;
wire \the_processor_cpu_nios2_ocimem|MonDReg[17]~q ;
wire \the_processor_cpu_nios2_ocimem|processor_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[5] ;
wire \the_processor_cpu_nios2_ocimem|processor_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[21] ;
wire \the_processor_cpu_nios2_ocimem|processor_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[13] ;
wire \the_processor_cpu_nios2_ocimem|processor_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[29] ;
wire \the_processor_cpu_nios2_ocimem|processor_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[4] ;
wire \the_processor_cpu_nios2_ocimem|processor_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[12] ;
wire \the_processor_cpu_nios2_ocimem|processor_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[28] ;
wire \the_processor_cpu_nios2_ocimem|processor_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[6] ;
wire \the_processor_cpu_nios2_ocimem|processor_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[22] ;
wire \the_processor_cpu_nios2_ocimem|processor_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[14] ;
wire \the_processor_cpu_nios2_ocimem|processor_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[30] ;
wire \the_processor_cpu_nios2_ocimem|processor_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[7] ;
wire \the_processor_cpu_nios2_ocimem|processor_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[23] ;
wire \the_processor_cpu_nios2_ocimem|processor_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[15] ;
wire \the_processor_cpu_nios2_ocimem|processor_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[31] ;
wire \the_processor_cpu_nios2_ocimem|processor_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[11] ;
wire \the_processor_cpu_nios2_ocimem|processor_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[27] ;
wire \the_processor_cpu_nios2_ocimem|processor_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[10] ;
wire \the_processor_cpu_nios2_ocimem|processor_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[26] ;
wire \the_processor_cpu_nios2_ocimem|processor_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[25] ;
wire \the_processor_cpu_nios2_ocimem|processor_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[9] ;
wire \the_processor_cpu_nios2_ocimem|processor_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[3] ;
wire \the_processor_cpu_nios2_ocimem|processor_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[18] ;
wire \the_processor_cpu_nios2_ocimem|processor_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[17] ;
wire \the_processor_cpu_nios2_oci_break|break_readreg[24]~q ;
wire \the_processor_cpu_nios2_ocimem|MonDReg[24]~q ;
wire \the_processor_cpu_nios2_oci_break|break_readreg[4]~q ;
wire \the_processor_cpu_nios2_oci_break|break_readreg[26]~q ;
wire \the_processor_cpu_nios2_ocimem|MonDReg[26]~q ;
wire \the_processor_cpu_nios2_oci_break|break_readreg[25]~q ;
wire \the_processor_cpu_nios2_ocimem|MonDReg[25]~q ;
wire \the_processor_cpu_nios2_oci_break|break_readreg[27]~q ;
wire \the_processor_cpu_nios2_ocimem|MonDReg[27]~q ;
wire \the_processor_cpu_nios2_oci_break|break_readreg[22]~q ;
wire \the_processor_cpu_nios2_ocimem|MonDReg[22]~q ;
wire \the_processor_cpu_nios2_ocimem|MonDReg[13]~q ;
wire \the_processor_cpu_nios2_ocimem|MonDReg[28]~q ;
wire \the_processor_cpu_nios2_ocimem|MonDReg[6]~q ;
wire \the_processor_cpu_nios2_ocimem|MonDReg[14]~q ;
wire \the_processor_cpu_nios2_ocimem|MonDReg[30]~q ;
wire \the_processor_cpu_nios2_ocimem|MonDReg[7]~q ;
wire \the_processor_cpu_nios2_ocimem|MonDReg[23]~q ;
wire \the_processor_cpu_nios2_ocimem|MonDReg[31]~q ;
wire \the_processor_cpu_nios2_ocimem|MonDReg[11]~q ;
wire \the_processor_cpu_nios2_ocimem|MonDReg[10]~q ;
wire \the_processor_cpu_nios2_ocimem|MonDReg[9]~q ;
wire \the_processor_cpu_nios2_oci_break|break_readreg[5]~q ;
wire \the_processor_cpu_nios2_oci_break|break_readreg[28]~q ;
wire \the_processor_cpu_nios2_oci_break|break_readreg[29]~q ;
wire \the_processor_cpu_nios2_oci_break|break_readreg[30]~q ;
wire \the_processor_cpu_nios2_oci_break|break_readreg[31]~q ;
wire \the_processor_cpu_nios2_oci_break|break_readreg[23]~q ;
wire \the_processor_cpu_nios2_oci_break|break_readreg[6]~q ;
wire \the_processor_cpu_nios2_oci_break|break_readreg[15]~q ;
wire \the_processor_cpu_nios2_oci_break|break_readreg[7]~q ;
wire \the_processor_cpu_nios2_oci_break|break_readreg[10]~q ;
wire \the_processor_cpu_nios2_oci_break|break_readreg[14]~q ;
wire \the_processor_cpu_nios2_oci_break|break_readreg[8]~q ;
wire \the_processor_cpu_nios2_oci_break|break_readreg[9]~q ;
wire \the_processor_cpu_nios2_oci_break|break_readreg[13]~q ;
wire \the_processor_cpu_nios2_oci_break|break_readreg[12]~q ;
wire \the_processor_cpu_nios2_oci_break|break_readreg[11]~q ;
wire \the_processor_cpu_nios2_ocimem|MonDReg[0]~q ;
wire \write~q ;
wire \read~q ;
wire \the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[34]~q ;
wire \the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[35]~q ;
wire \the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|ir[1]~q ;
wire \the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|ir[0]~q ;
wire \the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|enable_action_strobe~q ;
wire \the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|take_action_ocimem_a~0_combout ;
wire \the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|take_action_ocimem_a~1_combout ;
wire \the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|take_action_ocimem_a~combout ;
wire \the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[21]~q ;
wire \the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[20]~q ;
wire \the_processor_cpu_nios2_oci_debug|monitor_ready~q ;
wire \the_processor_cpu_nios2_ocimem|MonDReg[1]~q ;
wire \the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[0]~q ;
wire \the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[36]~q ;
wire \the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[37]~q ;
wire \the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[3]~q ;
wire \write~0_combout ;
wire \write~1_combout ;
wire \write~2_combout ;
wire \the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[17]~q ;
wire \read~0_combout ;
wire \writedata[3]~q ;
wire \address[0]~q ;
wire \address[3]~q ;
wire \address[2]~q ;
wire \address[1]~q ;
wire \address[7]~q ;
wire \address[6]~q ;
wire \address[5]~q ;
wire \address[4]~q ;
wire \the_processor_cpu_nios2_avalon_reg|Equal0~1_combout ;
wire \debugaccess~q ;
wire \the_processor_cpu_nios2_avalon_reg|take_action_ocireg~0_combout ;
wire \the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[19]~q ;
wire \the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[18]~q ;
wire \the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[25]~q ;
wire \writedata[0]~q ;
wire \the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[1]~q ;
wire \the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[4]~q ;
wire \the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[27]~q ;
wire \the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[26]~q ;
wire \the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[28]~q ;
wire \byteenable[0]~q ;
wire \the_processor_cpu_nios2_oci_debug|monitor_error~q ;
wire \writedata[16]~q ;
wire \the_processor_cpu_nios2_avalon_reg|Equal1~0_combout ;
wire \the_processor_cpu_nios2_ocimem|MonDReg[3]~q ;
wire \the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[2]~q ;
wire \the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[5]~q ;
wire \writedata[1]~q ;
wire \the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[29]~q ;
wire \the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[30]~q ;
wire \the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[31]~q ;
wire \the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[32]~q ;
wire \the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[33]~q ;
wire \the_processor_cpu_nios2_avalon_reg|oci_ienable[0]~q ;
wire \the_processor_cpu_nios2_avalon_reg|oci_reg_readdata~0_combout ;
wire \the_processor_cpu_nios2_avalon_reg|oci_reg_readdata~1_combout ;
wire \the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[23]~q ;
wire \the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[22]~q ;
wire \the_processor_cpu_nios2_ocimem|MonDReg[18]~q ;
wire \the_processor_cpu_nios2_oci_debug|monitor_go~q ;
wire \the_processor_cpu_nios2_avalon_reg|oci_reg_readdata[1]~2_combout ;
wire \the_processor_cpu_nios2_ocimem|MonDReg[4]~q ;
wire \the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[6]~q ;
wire \writedata[2]~q ;
wire \byteenable[2]~q ;
wire \the_processor_cpu_nios2_ocimem|MonDReg[8]~q ;
wire \writedata[8]~q ;
wire \byteenable[1]~q ;
wire \writedata[24]~q ;
wire \byteenable[3]~q ;
wire \the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[16]~q ;
wire \the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[24]~q ;
wire \writedata[20]~q ;
wire \writedata[19]~q ;
wire \the_processor_cpu_nios2_ocimem|MonDReg[5]~q ;
wire \writedata[5]~q ;
wire \writedata[21]~q ;
wire \writedata[13]~q ;
wire \the_processor_cpu_nios2_ocimem|MonDReg[29]~q ;
wire \writedata[29]~q ;
wire \writedata[4]~q ;
wire \the_processor_cpu_nios2_ocimem|MonDReg[12]~q ;
wire \writedata[12]~q ;
wire \writedata[28]~q ;
wire \writedata[6]~q ;
wire \writedata[22]~q ;
wire \writedata[14]~q ;
wire \writedata[30]~q ;
wire \writedata[7]~q ;
wire \writedata[23]~q ;
wire \the_processor_cpu_nios2_ocimem|MonDReg[15]~q ;
wire \writedata[15]~q ;
wire \writedata[31]~q ;
wire \writedata[11]~q ;
wire \writedata[27]~q ;
wire \writedata[10]~q ;
wire \writedata[26]~q ;
wire \writedata[25]~q ;
wire \writedata[9]~q ;
wire \writedata[18]~q ;
wire \writedata[17]~q ;
wire \the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[7]~q ;
wire \the_processor_cpu_nios2_oci_debug|resetlatch~q ;
wire \the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[11]~q ;
wire \the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[8]~q ;
wire \the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[15]~q ;
wire \the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[9]~q ;
wire \the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[10]~q ;
wire \the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[14]~q ;
wire \the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[13]~q ;
wire \the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[12]~q ;
wire \readdata~0_combout ;
wire \address[8]~q ;
wire \readdata~1_combout ;
wire \readdata~2_combout ;


processor_processor_cpu_nios2_oci_debug the_processor_cpu_nios2_oci_debug(
	.r_sync_rst(r_sync_rst),
	.jtag_break1(jtag_break),
	.jdo_34(\the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[34]~q ),
	.jdo_35(\the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[35]~q ),
	.take_action_ocimem_a(\the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|take_action_ocimem_a~0_combout ),
	.take_action_ocimem_a1(\the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|take_action_ocimem_a~combout ),
	.jdo_21(\the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[21]~q ),
	.jdo_20(\the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[20]~q ),
	.monitor_ready1(\the_processor_cpu_nios2_oci_debug|monitor_ready~q ),
	.take_action_ocireg(\the_processor_cpu_nios2_avalon_reg|take_action_ocireg~0_combout ),
	.jdo_19(\the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[19]~q ),
	.jdo_18(\the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[18]~q ),
	.jdo_25(\the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[25]~q ),
	.writedata_0(\writedata[0]~q ),
	.monitor_error1(\the_processor_cpu_nios2_oci_debug|monitor_error~q ),
	.writedata_1(\writedata[1]~q ),
	.jdo_23(\the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[23]~q ),
	.monitor_go1(\the_processor_cpu_nios2_oci_debug|monitor_go~q ),
	.jdo_24(\the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[24]~q ),
	.resetlatch1(\the_processor_cpu_nios2_oci_debug|resetlatch~q ),
	.state_1(state_1),
	.clk_clk(clk_clk));

processor_processor_cpu_nios2_oci_break the_processor_cpu_nios2_oci_break(
	.break_readreg_0(\the_processor_cpu_nios2_oci_break|break_readreg[0]~q ),
	.break_readreg_1(\the_processor_cpu_nios2_oci_break|break_readreg[1]~q ),
	.break_readreg_2(\the_processor_cpu_nios2_oci_break|break_readreg[2]~q ),
	.break_readreg_20(\the_processor_cpu_nios2_oci_break|break_readreg[20]~q ),
	.break_readreg_19(\the_processor_cpu_nios2_oci_break|break_readreg[19]~q ),
	.break_readreg_3(\the_processor_cpu_nios2_oci_break|break_readreg[3]~q ),
	.break_readreg_16(\the_processor_cpu_nios2_oci_break|break_readreg[16]~q ),
	.break_readreg_21(\the_processor_cpu_nios2_oci_break|break_readreg[21]~q ),
	.break_readreg_18(\the_processor_cpu_nios2_oci_break|break_readreg[18]~q ),
	.break_readreg_17(\the_processor_cpu_nios2_oci_break|break_readreg[17]~q ),
	.break_readreg_24(\the_processor_cpu_nios2_oci_break|break_readreg[24]~q ),
	.break_readreg_4(\the_processor_cpu_nios2_oci_break|break_readreg[4]~q ),
	.break_readreg_26(\the_processor_cpu_nios2_oci_break|break_readreg[26]~q ),
	.break_readreg_25(\the_processor_cpu_nios2_oci_break|break_readreg[25]~q ),
	.break_readreg_27(\the_processor_cpu_nios2_oci_break|break_readreg[27]~q ),
	.break_readreg_22(\the_processor_cpu_nios2_oci_break|break_readreg[22]~q ),
	.break_readreg_5(\the_processor_cpu_nios2_oci_break|break_readreg[5]~q ),
	.break_readreg_28(\the_processor_cpu_nios2_oci_break|break_readreg[28]~q ),
	.break_readreg_29(\the_processor_cpu_nios2_oci_break|break_readreg[29]~q ),
	.break_readreg_30(\the_processor_cpu_nios2_oci_break|break_readreg[30]~q ),
	.break_readreg_31(\the_processor_cpu_nios2_oci_break|break_readreg[31]~q ),
	.break_readreg_23(\the_processor_cpu_nios2_oci_break|break_readreg[23]~q ),
	.break_readreg_6(\the_processor_cpu_nios2_oci_break|break_readreg[6]~q ),
	.break_readreg_15(\the_processor_cpu_nios2_oci_break|break_readreg[15]~q ),
	.break_readreg_7(\the_processor_cpu_nios2_oci_break|break_readreg[7]~q ),
	.break_readreg_10(\the_processor_cpu_nios2_oci_break|break_readreg[10]~q ),
	.break_readreg_14(\the_processor_cpu_nios2_oci_break|break_readreg[14]~q ),
	.break_readreg_8(\the_processor_cpu_nios2_oci_break|break_readreg[8]~q ),
	.break_readreg_9(\the_processor_cpu_nios2_oci_break|break_readreg[9]~q ),
	.break_readreg_13(\the_processor_cpu_nios2_oci_break|break_readreg[13]~q ),
	.break_readreg_12(\the_processor_cpu_nios2_oci_break|break_readreg[12]~q ),
	.break_readreg_11(\the_processor_cpu_nios2_oci_break|break_readreg[11]~q ),
	.ir_1(\the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|ir[1]~q ),
	.ir_0(\the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|ir[0]~q ),
	.enable_action_strobe(\the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|enable_action_strobe~q ),
	.jdo_21(\the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[21]~q ),
	.jdo_20(\the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[20]~q ),
	.jdo_0(\the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[0]~q ),
	.jdo_36(\the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[36]~q ),
	.jdo_37(\the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[37]~q ),
	.jdo_3(\the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[3]~q ),
	.jdo_17(\the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[17]~q ),
	.jdo_19(\the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[19]~q ),
	.jdo_18(\the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[18]~q ),
	.jdo_25(\the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[25]~q ),
	.jdo_1(\the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[1]~q ),
	.jdo_4(\the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[4]~q ),
	.jdo_27(\the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[27]~q ),
	.jdo_26(\the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[26]~q ),
	.jdo_28(\the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[28]~q ),
	.jdo_2(\the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[2]~q ),
	.jdo_5(\the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[5]~q ),
	.jdo_29(\the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[29]~q ),
	.jdo_30(\the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[30]~q ),
	.jdo_31(\the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[31]~q ),
	.jdo_23(\the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[23]~q ),
	.jdo_22(\the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[22]~q ),
	.jdo_6(\the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[6]~q ),
	.jdo_16(\the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[16]~q ),
	.jdo_24(\the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[24]~q ),
	.jdo_7(\the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[7]~q ),
	.jdo_11(\the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[11]~q ),
	.jdo_8(\the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[8]~q ),
	.jdo_15(\the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[15]~q ),
	.jdo_9(\the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[9]~q ),
	.jdo_10(\the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[10]~q ),
	.jdo_14(\the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[14]~q ),
	.jdo_13(\the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[13]~q ),
	.jdo_12(\the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[12]~q ),
	.clk_clk(clk_clk));

processor_processor_cpu_nios2_avalon_reg the_processor_cpu_nios2_avalon_reg(
	.r_sync_rst(r_sync_rst),
	.write(\write~q ),
	.address_8(\address[8]~q ),
	.oci_single_step_mode1(oci_single_step_mode),
	.monitor_ready(\the_processor_cpu_nios2_oci_debug|monitor_ready~q ),
	.writedata_3(\writedata[3]~q ),
	.address_0(\address[0]~q ),
	.address_3(\address[3]~q ),
	.address_2(\address[2]~q ),
	.address_1(\address[1]~q ),
	.address_7(\address[7]~q ),
	.address_6(\address[6]~q ),
	.address_5(\address[5]~q ),
	.address_4(\address[4]~q ),
	.Equal0(\the_processor_cpu_nios2_avalon_reg|Equal0~1_combout ),
	.debugaccess(\debugaccess~q ),
	.take_action_ocireg(\the_processor_cpu_nios2_avalon_reg|take_action_ocireg~0_combout ),
	.oci_ienable_16(oci_ienable_16),
	.oci_ienable_1(oci_ienable_1),
	.writedata_16(\writedata[16]~q ),
	.Equal1(\the_processor_cpu_nios2_avalon_reg|Equal1~0_combout ),
	.writedata_1(\writedata[1]~q ),
	.oci_ienable_0(\the_processor_cpu_nios2_avalon_reg|oci_ienable[0]~q ),
	.oci_reg_readdata(\the_processor_cpu_nios2_avalon_reg|oci_reg_readdata~0_combout ),
	.oci_reg_readdata1(\the_processor_cpu_nios2_avalon_reg|oci_reg_readdata~1_combout ),
	.oci_reg_readdata_1(\the_processor_cpu_nios2_avalon_reg|oci_reg_readdata[1]~2_combout ),
	.clk_clk(clk_clk));

processor_processor_cpu_nios2_ocimem the_processor_cpu_nios2_ocimem(
	.q_a_0(\the_processor_cpu_nios2_ocimem|processor_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[0] ),
	.MonDReg_2(\the_processor_cpu_nios2_ocimem|MonDReg[2]~q ),
	.q_a_1(\the_processor_cpu_nios2_ocimem|processor_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[1] ),
	.MonDReg_20(\the_processor_cpu_nios2_ocimem|MonDReg[20]~q ),
	.MonDReg_19(\the_processor_cpu_nios2_ocimem|MonDReg[19]~q ),
	.q_a_2(\the_processor_cpu_nios2_ocimem|processor_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[2] ),
	.q_a_16(\the_processor_cpu_nios2_ocimem|processor_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[16] ),
	.q_a_8(\the_processor_cpu_nios2_ocimem|processor_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[8] ),
	.q_a_24(\the_processor_cpu_nios2_ocimem|processor_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[24] ),
	.MonDReg_16(\the_processor_cpu_nios2_ocimem|MonDReg[16]~q ),
	.MonDReg_21(\the_processor_cpu_nios2_ocimem|MonDReg[21]~q ),
	.q_a_20(\the_processor_cpu_nios2_ocimem|processor_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[20] ),
	.q_a_19(\the_processor_cpu_nios2_ocimem|processor_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[19] ),
	.MonDReg_17(\the_processor_cpu_nios2_ocimem|MonDReg[17]~q ),
	.q_a_5(\the_processor_cpu_nios2_ocimem|processor_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[5] ),
	.q_a_21(\the_processor_cpu_nios2_ocimem|processor_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[21] ),
	.q_a_13(\the_processor_cpu_nios2_ocimem|processor_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[13] ),
	.q_a_29(\the_processor_cpu_nios2_ocimem|processor_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[29] ),
	.q_a_4(\the_processor_cpu_nios2_ocimem|processor_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[4] ),
	.q_a_12(\the_processor_cpu_nios2_ocimem|processor_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[12] ),
	.q_a_28(\the_processor_cpu_nios2_ocimem|processor_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[28] ),
	.q_a_6(\the_processor_cpu_nios2_ocimem|processor_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[6] ),
	.q_a_22(\the_processor_cpu_nios2_ocimem|processor_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[22] ),
	.q_a_14(\the_processor_cpu_nios2_ocimem|processor_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[14] ),
	.q_a_30(\the_processor_cpu_nios2_ocimem|processor_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[30] ),
	.q_a_7(\the_processor_cpu_nios2_ocimem|processor_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[7] ),
	.q_a_23(\the_processor_cpu_nios2_ocimem|processor_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[23] ),
	.q_a_15(\the_processor_cpu_nios2_ocimem|processor_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[15] ),
	.q_a_31(\the_processor_cpu_nios2_ocimem|processor_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[31] ),
	.q_a_11(\the_processor_cpu_nios2_ocimem|processor_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[11] ),
	.q_a_27(\the_processor_cpu_nios2_ocimem|processor_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[27] ),
	.q_a_10(\the_processor_cpu_nios2_ocimem|processor_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[10] ),
	.q_a_26(\the_processor_cpu_nios2_ocimem|processor_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[26] ),
	.q_a_25(\the_processor_cpu_nios2_ocimem|processor_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[25] ),
	.q_a_9(\the_processor_cpu_nios2_ocimem|processor_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[9] ),
	.q_a_3(\the_processor_cpu_nios2_ocimem|processor_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[3] ),
	.q_a_18(\the_processor_cpu_nios2_ocimem|processor_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[18] ),
	.q_a_17(\the_processor_cpu_nios2_ocimem|processor_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[17] ),
	.MonDReg_24(\the_processor_cpu_nios2_ocimem|MonDReg[24]~q ),
	.MonDReg_26(\the_processor_cpu_nios2_ocimem|MonDReg[26]~q ),
	.MonDReg_25(\the_processor_cpu_nios2_ocimem|MonDReg[25]~q ),
	.MonDReg_27(\the_processor_cpu_nios2_ocimem|MonDReg[27]~q ),
	.MonDReg_22(\the_processor_cpu_nios2_ocimem|MonDReg[22]~q ),
	.MonDReg_13(\the_processor_cpu_nios2_ocimem|MonDReg[13]~q ),
	.MonDReg_28(\the_processor_cpu_nios2_ocimem|MonDReg[28]~q ),
	.MonDReg_6(\the_processor_cpu_nios2_ocimem|MonDReg[6]~q ),
	.MonDReg_14(\the_processor_cpu_nios2_ocimem|MonDReg[14]~q ),
	.MonDReg_30(\the_processor_cpu_nios2_ocimem|MonDReg[30]~q ),
	.MonDReg_7(\the_processor_cpu_nios2_ocimem|MonDReg[7]~q ),
	.MonDReg_23(\the_processor_cpu_nios2_ocimem|MonDReg[23]~q ),
	.MonDReg_31(\the_processor_cpu_nios2_ocimem|MonDReg[31]~q ),
	.MonDReg_11(\the_processor_cpu_nios2_ocimem|MonDReg[11]~q ),
	.MonDReg_10(\the_processor_cpu_nios2_ocimem|MonDReg[10]~q ),
	.MonDReg_9(\the_processor_cpu_nios2_ocimem|MonDReg[9]~q ),
	.waitrequest1(waitrequest),
	.MonDReg_0(\the_processor_cpu_nios2_ocimem|MonDReg[0]~q ),
	.write(\write~q ),
	.address_8(\address[8]~q ),
	.read(\read~q ),
	.jdo_34(\the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[34]~q ),
	.jdo_35(\the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[35]~q ),
	.take_action_ocimem_a(\the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|take_action_ocimem_a~0_combout ),
	.take_no_action_ocimem_a(\the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|take_action_ocimem_a~1_combout ),
	.take_action_ocimem_a1(\the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|take_action_ocimem_a~combout ),
	.jdo_21(\the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[21]~q ),
	.jdo_20(\the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[20]~q ),
	.MonDReg_1(\the_processor_cpu_nios2_ocimem|MonDReg[1]~q ),
	.jdo_3(\the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[3]~q ),
	.jdo_17(\the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[17]~q ),
	.writedata_3(\writedata[3]~q ),
	.address_0(\address[0]~q ),
	.address_3(\address[3]~q ),
	.address_2(\address[2]~q ),
	.address_1(\address[1]~q ),
	.address_7(\address[7]~q ),
	.address_6(\address[6]~q ),
	.address_5(\address[5]~q ),
	.address_4(\address[4]~q ),
	.debugaccess(\debugaccess~q ),
	.jdo_19(\the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[19]~q ),
	.jdo_18(\the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[18]~q ),
	.jdo_25(\the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[25]~q ),
	.writedata_0(\writedata[0]~q ),
	.jdo_4(\the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[4]~q ),
	.jdo_27(\the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[27]~q ),
	.jdo_26(\the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[26]~q ),
	.jdo_28(\the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[28]~q ),
	.r_early_rst(r_early_rst),
	.byteenable_0(\byteenable[0]~q ),
	.writedata_16(\writedata[16]~q ),
	.MonDReg_3(\the_processor_cpu_nios2_ocimem|MonDReg[3]~q ),
	.jdo_5(\the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[5]~q ),
	.writedata_1(\writedata[1]~q ),
	.jdo_29(\the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[29]~q ),
	.jdo_30(\the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[30]~q ),
	.jdo_31(\the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[31]~q ),
	.jdo_32(\the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[32]~q ),
	.jdo_33(\the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[33]~q ),
	.jdo_23(\the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[23]~q ),
	.jdo_22(\the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[22]~q ),
	.MonDReg_18(\the_processor_cpu_nios2_ocimem|MonDReg[18]~q ),
	.MonDReg_4(\the_processor_cpu_nios2_ocimem|MonDReg[4]~q ),
	.jdo_6(\the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[6]~q ),
	.writedata_2(\writedata[2]~q ),
	.byteenable_2(\byteenable[2]~q ),
	.MonDReg_8(\the_processor_cpu_nios2_ocimem|MonDReg[8]~q ),
	.writedata_8(\writedata[8]~q ),
	.byteenable_1(\byteenable[1]~q ),
	.writedata_24(\writedata[24]~q ),
	.byteenable_3(\byteenable[3]~q ),
	.jdo_16(\the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[16]~q ),
	.jdo_24(\the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[24]~q ),
	.writedata_20(\writedata[20]~q ),
	.writedata_19(\writedata[19]~q ),
	.MonDReg_5(\the_processor_cpu_nios2_ocimem|MonDReg[5]~q ),
	.writedata_5(\writedata[5]~q ),
	.writedata_21(\writedata[21]~q ),
	.writedata_13(\writedata[13]~q ),
	.MonDReg_29(\the_processor_cpu_nios2_ocimem|MonDReg[29]~q ),
	.writedata_29(\writedata[29]~q ),
	.writedata_4(\writedata[4]~q ),
	.MonDReg_12(\the_processor_cpu_nios2_ocimem|MonDReg[12]~q ),
	.writedata_12(\writedata[12]~q ),
	.writedata_28(\writedata[28]~q ),
	.writedata_6(\writedata[6]~q ),
	.writedata_22(\writedata[22]~q ),
	.writedata_14(\writedata[14]~q ),
	.writedata_30(\writedata[30]~q ),
	.writedata_7(\writedata[7]~q ),
	.writedata_23(\writedata[23]~q ),
	.MonDReg_15(\the_processor_cpu_nios2_ocimem|MonDReg[15]~q ),
	.writedata_15(\writedata[15]~q ),
	.writedata_31(\writedata[31]~q ),
	.writedata_11(\writedata[11]~q ),
	.writedata_27(\writedata[27]~q ),
	.writedata_10(\writedata[10]~q ),
	.writedata_26(\writedata[26]~q ),
	.writedata_25(\writedata[25]~q ),
	.writedata_9(\writedata[9]~q ),
	.writedata_18(\writedata[18]~q ),
	.writedata_17(\writedata[17]~q ),
	.jdo_7(\the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[7]~q ),
	.jdo_11(\the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[11]~q ),
	.jdo_8(\the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[8]~q ),
	.jdo_15(\the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[15]~q ),
	.jdo_9(\the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[9]~q ),
	.jdo_10(\the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[10]~q ),
	.jdo_14(\the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[14]~q ),
	.jdo_13(\the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[13]~q ),
	.jdo_12(\the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[12]~q ),
	.clk_clk(clk_clk));

processor_processor_cpu_jtag_debug_module_wrapper the_processor_cpu_jtag_debug_module_wrapper(
	.break_readreg_0(\the_processor_cpu_nios2_oci_break|break_readreg[0]~q ),
	.break_readreg_1(\the_processor_cpu_nios2_oci_break|break_readreg[1]~q ),
	.break_readreg_2(\the_processor_cpu_nios2_oci_break|break_readreg[2]~q ),
	.MonDReg_2(\the_processor_cpu_nios2_ocimem|MonDReg[2]~q ),
	.break_readreg_20(\the_processor_cpu_nios2_oci_break|break_readreg[20]~q ),
	.MonDReg_20(\the_processor_cpu_nios2_ocimem|MonDReg[20]~q ),
	.break_readreg_19(\the_processor_cpu_nios2_oci_break|break_readreg[19]~q ),
	.MonDReg_19(\the_processor_cpu_nios2_ocimem|MonDReg[19]~q ),
	.break_readreg_3(\the_processor_cpu_nios2_oci_break|break_readreg[3]~q ),
	.break_readreg_16(\the_processor_cpu_nios2_oci_break|break_readreg[16]~q ),
	.MonDReg_16(\the_processor_cpu_nios2_ocimem|MonDReg[16]~q ),
	.break_readreg_21(\the_processor_cpu_nios2_oci_break|break_readreg[21]~q ),
	.MonDReg_21(\the_processor_cpu_nios2_ocimem|MonDReg[21]~q ),
	.break_readreg_18(\the_processor_cpu_nios2_oci_break|break_readreg[18]~q ),
	.break_readreg_17(\the_processor_cpu_nios2_oci_break|break_readreg[17]~q ),
	.MonDReg_17(\the_processor_cpu_nios2_ocimem|MonDReg[17]~q ),
	.break_readreg_24(\the_processor_cpu_nios2_oci_break|break_readreg[24]~q ),
	.MonDReg_24(\the_processor_cpu_nios2_ocimem|MonDReg[24]~q ),
	.break_readreg_4(\the_processor_cpu_nios2_oci_break|break_readreg[4]~q ),
	.break_readreg_26(\the_processor_cpu_nios2_oci_break|break_readreg[26]~q ),
	.MonDReg_26(\the_processor_cpu_nios2_ocimem|MonDReg[26]~q ),
	.break_readreg_25(\the_processor_cpu_nios2_oci_break|break_readreg[25]~q ),
	.MonDReg_25(\the_processor_cpu_nios2_ocimem|MonDReg[25]~q ),
	.break_readreg_27(\the_processor_cpu_nios2_oci_break|break_readreg[27]~q ),
	.MonDReg_27(\the_processor_cpu_nios2_ocimem|MonDReg[27]~q ),
	.break_readreg_22(\the_processor_cpu_nios2_oci_break|break_readreg[22]~q ),
	.MonDReg_22(\the_processor_cpu_nios2_ocimem|MonDReg[22]~q ),
	.MonDReg_13(\the_processor_cpu_nios2_ocimem|MonDReg[13]~q ),
	.MonDReg_28(\the_processor_cpu_nios2_ocimem|MonDReg[28]~q ),
	.MonDReg_6(\the_processor_cpu_nios2_ocimem|MonDReg[6]~q ),
	.MonDReg_14(\the_processor_cpu_nios2_ocimem|MonDReg[14]~q ),
	.MonDReg_30(\the_processor_cpu_nios2_ocimem|MonDReg[30]~q ),
	.MonDReg_7(\the_processor_cpu_nios2_ocimem|MonDReg[7]~q ),
	.MonDReg_23(\the_processor_cpu_nios2_ocimem|MonDReg[23]~q ),
	.MonDReg_31(\the_processor_cpu_nios2_ocimem|MonDReg[31]~q ),
	.MonDReg_11(\the_processor_cpu_nios2_ocimem|MonDReg[11]~q ),
	.MonDReg_10(\the_processor_cpu_nios2_ocimem|MonDReg[10]~q ),
	.MonDReg_9(\the_processor_cpu_nios2_ocimem|MonDReg[9]~q ),
	.break_readreg_5(\the_processor_cpu_nios2_oci_break|break_readreg[5]~q ),
	.break_readreg_28(\the_processor_cpu_nios2_oci_break|break_readreg[28]~q ),
	.break_readreg_29(\the_processor_cpu_nios2_oci_break|break_readreg[29]~q ),
	.break_readreg_30(\the_processor_cpu_nios2_oci_break|break_readreg[30]~q ),
	.break_readreg_31(\the_processor_cpu_nios2_oci_break|break_readreg[31]~q ),
	.break_readreg_23(\the_processor_cpu_nios2_oci_break|break_readreg[23]~q ),
	.break_readreg_6(\the_processor_cpu_nios2_oci_break|break_readreg[6]~q ),
	.break_readreg_15(\the_processor_cpu_nios2_oci_break|break_readreg[15]~q ),
	.break_readreg_7(\the_processor_cpu_nios2_oci_break|break_readreg[7]~q ),
	.break_readreg_10(\the_processor_cpu_nios2_oci_break|break_readreg[10]~q ),
	.break_readreg_14(\the_processor_cpu_nios2_oci_break|break_readreg[14]~q ),
	.break_readreg_8(\the_processor_cpu_nios2_oci_break|break_readreg[8]~q ),
	.break_readreg_9(\the_processor_cpu_nios2_oci_break|break_readreg[9]~q ),
	.break_readreg_13(\the_processor_cpu_nios2_oci_break|break_readreg[13]~q ),
	.break_readreg_12(\the_processor_cpu_nios2_oci_break|break_readreg[12]~q ),
	.break_readreg_11(\the_processor_cpu_nios2_oci_break|break_readreg[11]~q ),
	.sr_0(sr_0),
	.ir_out_0(ir_out_0),
	.ir_out_1(ir_out_1),
	.hbreak_enabled(hbreak_enabled),
	.MonDReg_0(\the_processor_cpu_nios2_ocimem|MonDReg[0]~q ),
	.jdo_34(\the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[34]~q ),
	.jdo_35(\the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[35]~q ),
	.ir_1(\the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|ir[1]~q ),
	.ir_0(\the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|ir[0]~q ),
	.enable_action_strobe(\the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|enable_action_strobe~q ),
	.take_action_ocimem_a(\the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|take_action_ocimem_a~0_combout ),
	.take_action_ocimem_a1(\the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|take_action_ocimem_a~1_combout ),
	.take_action_ocimem_a2(\the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|take_action_ocimem_a~combout ),
	.jdo_21(\the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[21]~q ),
	.jdo_20(\the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[20]~q ),
	.monitor_ready(\the_processor_cpu_nios2_oci_debug|monitor_ready~q ),
	.MonDReg_1(\the_processor_cpu_nios2_ocimem|MonDReg[1]~q ),
	.jdo_0(\the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[0]~q ),
	.jdo_36(\the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[36]~q ),
	.jdo_37(\the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[37]~q ),
	.jdo_3(\the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[3]~q ),
	.jdo_17(\the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[17]~q ),
	.jdo_19(\the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[19]~q ),
	.jdo_18(\the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[18]~q ),
	.jdo_25(\the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[25]~q ),
	.jdo_1(\the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[1]~q ),
	.jdo_4(\the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[4]~q ),
	.jdo_27(\the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[27]~q ),
	.jdo_26(\the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[26]~q ),
	.jdo_28(\the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[28]~q ),
	.monitor_error(\the_processor_cpu_nios2_oci_debug|monitor_error~q ),
	.MonDReg_3(\the_processor_cpu_nios2_ocimem|MonDReg[3]~q ),
	.jdo_2(\the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[2]~q ),
	.jdo_5(\the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[5]~q ),
	.jdo_29(\the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[29]~q ),
	.jdo_30(\the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[30]~q ),
	.jdo_31(\the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[31]~q ),
	.jdo_32(\the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[32]~q ),
	.jdo_33(\the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[33]~q ),
	.jdo_23(\the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[23]~q ),
	.jdo_22(\the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[22]~q ),
	.MonDReg_18(\the_processor_cpu_nios2_ocimem|MonDReg[18]~q ),
	.MonDReg_4(\the_processor_cpu_nios2_ocimem|MonDReg[4]~q ),
	.jdo_6(\the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[6]~q ),
	.MonDReg_8(\the_processor_cpu_nios2_ocimem|MonDReg[8]~q ),
	.jdo_16(\the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[16]~q ),
	.jdo_24(\the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[24]~q ),
	.MonDReg_5(\the_processor_cpu_nios2_ocimem|MonDReg[5]~q ),
	.MonDReg_29(\the_processor_cpu_nios2_ocimem|MonDReg[29]~q ),
	.MonDReg_12(\the_processor_cpu_nios2_ocimem|MonDReg[12]~q ),
	.MonDReg_15(\the_processor_cpu_nios2_ocimem|MonDReg[15]~q ),
	.jdo_7(\the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[7]~q ),
	.resetlatch(\the_processor_cpu_nios2_oci_debug|resetlatch~q ),
	.jdo_11(\the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[11]~q ),
	.jdo_8(\the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[8]~q ),
	.jdo_15(\the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[15]~q ),
	.jdo_9(\the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[9]~q ),
	.jdo_10(\the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[10]~q ),
	.jdo_14(\the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[14]~q ),
	.jdo_13(\the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[13]~q ),
	.jdo_12(\the_processor_cpu_jtag_debug_module_wrapper|the_processor_cpu_jtag_debug_module_sysclk|jdo[12]~q ),
	.altera_internal_jtag(altera_internal_jtag),
	.altera_internal_jtag1(altera_internal_jtag1),
	.state_4(state_4),
	.virtual_ir_scan_reg(virtual_ir_scan_reg),
	.state_3(state_3),
	.state_8(state_8),
	.splitter_nodes_receive_1_3(splitter_nodes_receive_1_3),
	.irf_reg_0_2(irf_reg_0_2),
	.irf_reg_1_2(irf_reg_1_2),
	.clk_clk(clk_clk));

dffeas write(
	.clk(clk_clk),
	.d(\write~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\write~q ),
	.prn(vcc));
defparam write.is_wysiwyg = "true";
defparam write.power_up = "low";

dffeas read(
	.clk(clk_clk),
	.d(\read~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\read~q ),
	.prn(vcc));
defparam read.is_wysiwyg = "true";
defparam read.power_up = "low";

cyclonev_lcell_comb \write~0 (
	.dataa(!d_write),
	.datab(!mem_used_1),
	.datac(!\write~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\write~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \write~0 .extended_lut = "off";
defparam \write~0 .lut_mask = 64'hFDFDFDFDFDFDFDFD;
defparam \write~0 .shared_arith = "off";

cyclonev_lcell_comb \write~1 (
	.dataa(!saved_grant_0),
	.datab(!src2_valid),
	.datac(!saved_grant_1),
	.datad(!src0_valid),
	.datae(!\write~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\write~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \write~1 .extended_lut = "off";
defparam \write~1 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \write~1 .shared_arith = "off";

cyclonev_lcell_comb \write~2 (
	.dataa(!waitrequest),
	.datab(!\write~q ),
	.datac(!\write~1_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\write~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \write~2 .extended_lut = "off";
defparam \write~2 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \write~2 .shared_arith = "off";

cyclonev_lcell_comb \read~0 (
	.dataa(!waitrequest),
	.datab(!mem_used_1),
	.datac(!rf_source_valid),
	.datad(!\read~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read~0 .extended_lut = "off";
defparam \read~0 .lut_mask = 64'hCF5FCF5FCF5FCF5F;
defparam \read~0 .shared_arith = "off";

dffeas \writedata[3] (
	.clk(clk_clk),
	.d(writedata_nxt[3]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[3]~q ),
	.prn(vcc));
defparam \writedata[3] .is_wysiwyg = "true";
defparam \writedata[3] .power_up = "low";

dffeas \address[0] (
	.clk(clk_clk),
	.d(address_nxt[0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\address[0]~q ),
	.prn(vcc));
defparam \address[0] .is_wysiwyg = "true";
defparam \address[0] .power_up = "low";

dffeas \address[3] (
	.clk(clk_clk),
	.d(address_nxt[3]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\address[3]~q ),
	.prn(vcc));
defparam \address[3] .is_wysiwyg = "true";
defparam \address[3] .power_up = "low";

dffeas \address[2] (
	.clk(clk_clk),
	.d(address_nxt[2]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\address[2]~q ),
	.prn(vcc));
defparam \address[2] .is_wysiwyg = "true";
defparam \address[2] .power_up = "low";

dffeas \address[1] (
	.clk(clk_clk),
	.d(address_nxt[1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\address[1]~q ),
	.prn(vcc));
defparam \address[1] .is_wysiwyg = "true";
defparam \address[1] .power_up = "low";

dffeas \address[7] (
	.clk(clk_clk),
	.d(address_nxt[7]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\address[7]~q ),
	.prn(vcc));
defparam \address[7] .is_wysiwyg = "true";
defparam \address[7] .power_up = "low";

dffeas \address[6] (
	.clk(clk_clk),
	.d(address_nxt[6]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\address[6]~q ),
	.prn(vcc));
defparam \address[6] .is_wysiwyg = "true";
defparam \address[6] .power_up = "low";

dffeas \address[5] (
	.clk(clk_clk),
	.d(address_nxt[5]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\address[5]~q ),
	.prn(vcc));
defparam \address[5] .is_wysiwyg = "true";
defparam \address[5] .power_up = "low";

dffeas \address[4] (
	.clk(clk_clk),
	.d(address_nxt[4]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\address[4]~q ),
	.prn(vcc));
defparam \address[4] .is_wysiwyg = "true";
defparam \address[4] .power_up = "low";

dffeas debugaccess(
	.clk(clk_clk),
	.d(debugaccess_nxt),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\debugaccess~q ),
	.prn(vcc));
defparam debugaccess.is_wysiwyg = "true";
defparam debugaccess.power_up = "low";

dffeas \writedata[0] (
	.clk(clk_clk),
	.d(writedata_nxt[0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[0]~q ),
	.prn(vcc));
defparam \writedata[0] .is_wysiwyg = "true";
defparam \writedata[0] .power_up = "low";

dffeas \byteenable[0] (
	.clk(clk_clk),
	.d(byteenable_nxt[0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\byteenable[0]~q ),
	.prn(vcc));
defparam \byteenable[0] .is_wysiwyg = "true";
defparam \byteenable[0] .power_up = "low";

dffeas \writedata[16] (
	.clk(clk_clk),
	.d(writedata_nxt[16]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[16]~q ),
	.prn(vcc));
defparam \writedata[16] .is_wysiwyg = "true";
defparam \writedata[16] .power_up = "low";

dffeas \writedata[1] (
	.clk(clk_clk),
	.d(writedata_nxt[1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[1]~q ),
	.prn(vcc));
defparam \writedata[1] .is_wysiwyg = "true";
defparam \writedata[1] .power_up = "low";

dffeas \writedata[2] (
	.clk(clk_clk),
	.d(writedata_nxt[2]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[2]~q ),
	.prn(vcc));
defparam \writedata[2] .is_wysiwyg = "true";
defparam \writedata[2] .power_up = "low";

dffeas \byteenable[2] (
	.clk(clk_clk),
	.d(byteenable_nxt[2]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\byteenable[2]~q ),
	.prn(vcc));
defparam \byteenable[2] .is_wysiwyg = "true";
defparam \byteenable[2] .power_up = "low";

dffeas \writedata[8] (
	.clk(clk_clk),
	.d(writedata_nxt[8]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[8]~q ),
	.prn(vcc));
defparam \writedata[8] .is_wysiwyg = "true";
defparam \writedata[8] .power_up = "low";

dffeas \byteenable[1] (
	.clk(clk_clk),
	.d(byteenable_nxt[1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\byteenable[1]~q ),
	.prn(vcc));
defparam \byteenable[1] .is_wysiwyg = "true";
defparam \byteenable[1] .power_up = "low";

dffeas \writedata[24] (
	.clk(clk_clk),
	.d(writedata_nxt[24]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[24]~q ),
	.prn(vcc));
defparam \writedata[24] .is_wysiwyg = "true";
defparam \writedata[24] .power_up = "low";

dffeas \byteenable[3] (
	.clk(clk_clk),
	.d(byteenable_nxt[3]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\byteenable[3]~q ),
	.prn(vcc));
defparam \byteenable[3] .is_wysiwyg = "true";
defparam \byteenable[3] .power_up = "low";

dffeas \writedata[20] (
	.clk(clk_clk),
	.d(writedata_nxt[20]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[20]~q ),
	.prn(vcc));
defparam \writedata[20] .is_wysiwyg = "true";
defparam \writedata[20] .power_up = "low";

dffeas \writedata[19] (
	.clk(clk_clk),
	.d(writedata_nxt[19]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[19]~q ),
	.prn(vcc));
defparam \writedata[19] .is_wysiwyg = "true";
defparam \writedata[19] .power_up = "low";

dffeas \writedata[5] (
	.clk(clk_clk),
	.d(writedata_nxt[5]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[5]~q ),
	.prn(vcc));
defparam \writedata[5] .is_wysiwyg = "true";
defparam \writedata[5] .power_up = "low";

dffeas \writedata[21] (
	.clk(clk_clk),
	.d(writedata_nxt[21]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[21]~q ),
	.prn(vcc));
defparam \writedata[21] .is_wysiwyg = "true";
defparam \writedata[21] .power_up = "low";

dffeas \writedata[13] (
	.clk(clk_clk),
	.d(writedata_nxt[13]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[13]~q ),
	.prn(vcc));
defparam \writedata[13] .is_wysiwyg = "true";
defparam \writedata[13] .power_up = "low";

dffeas \writedata[29] (
	.clk(clk_clk),
	.d(writedata_nxt[29]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[29]~q ),
	.prn(vcc));
defparam \writedata[29] .is_wysiwyg = "true";
defparam \writedata[29] .power_up = "low";

dffeas \writedata[4] (
	.clk(clk_clk),
	.d(writedata_nxt[4]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[4]~q ),
	.prn(vcc));
defparam \writedata[4] .is_wysiwyg = "true";
defparam \writedata[4] .power_up = "low";

dffeas \writedata[12] (
	.clk(clk_clk),
	.d(writedata_nxt[12]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[12]~q ),
	.prn(vcc));
defparam \writedata[12] .is_wysiwyg = "true";
defparam \writedata[12] .power_up = "low";

dffeas \writedata[28] (
	.clk(clk_clk),
	.d(writedata_nxt[28]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[28]~q ),
	.prn(vcc));
defparam \writedata[28] .is_wysiwyg = "true";
defparam \writedata[28] .power_up = "low";

dffeas \writedata[6] (
	.clk(clk_clk),
	.d(writedata_nxt[6]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[6]~q ),
	.prn(vcc));
defparam \writedata[6] .is_wysiwyg = "true";
defparam \writedata[6] .power_up = "low";

dffeas \writedata[22] (
	.clk(clk_clk),
	.d(writedata_nxt[22]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[22]~q ),
	.prn(vcc));
defparam \writedata[22] .is_wysiwyg = "true";
defparam \writedata[22] .power_up = "low";

dffeas \writedata[14] (
	.clk(clk_clk),
	.d(writedata_nxt[14]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[14]~q ),
	.prn(vcc));
defparam \writedata[14] .is_wysiwyg = "true";
defparam \writedata[14] .power_up = "low";

dffeas \writedata[30] (
	.clk(clk_clk),
	.d(writedata_nxt[30]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[30]~q ),
	.prn(vcc));
defparam \writedata[30] .is_wysiwyg = "true";
defparam \writedata[30] .power_up = "low";

dffeas \writedata[7] (
	.clk(clk_clk),
	.d(writedata_nxt[7]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[7]~q ),
	.prn(vcc));
defparam \writedata[7] .is_wysiwyg = "true";
defparam \writedata[7] .power_up = "low";

dffeas \writedata[23] (
	.clk(clk_clk),
	.d(writedata_nxt[23]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[23]~q ),
	.prn(vcc));
defparam \writedata[23] .is_wysiwyg = "true";
defparam \writedata[23] .power_up = "low";

dffeas \writedata[15] (
	.clk(clk_clk),
	.d(writedata_nxt[15]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[15]~q ),
	.prn(vcc));
defparam \writedata[15] .is_wysiwyg = "true";
defparam \writedata[15] .power_up = "low";

dffeas \writedata[31] (
	.clk(clk_clk),
	.d(writedata_nxt[31]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[31]~q ),
	.prn(vcc));
defparam \writedata[31] .is_wysiwyg = "true";
defparam \writedata[31] .power_up = "low";

dffeas \writedata[11] (
	.clk(clk_clk),
	.d(writedata_nxt[11]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[11]~q ),
	.prn(vcc));
defparam \writedata[11] .is_wysiwyg = "true";
defparam \writedata[11] .power_up = "low";

dffeas \writedata[27] (
	.clk(clk_clk),
	.d(writedata_nxt[27]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[27]~q ),
	.prn(vcc));
defparam \writedata[27] .is_wysiwyg = "true";
defparam \writedata[27] .power_up = "low";

dffeas \writedata[10] (
	.clk(clk_clk),
	.d(writedata_nxt[10]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[10]~q ),
	.prn(vcc));
defparam \writedata[10] .is_wysiwyg = "true";
defparam \writedata[10] .power_up = "low";

dffeas \writedata[26] (
	.clk(clk_clk),
	.d(writedata_nxt[26]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[26]~q ),
	.prn(vcc));
defparam \writedata[26] .is_wysiwyg = "true";
defparam \writedata[26] .power_up = "low";

dffeas \writedata[25] (
	.clk(clk_clk),
	.d(writedata_nxt[25]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[25]~q ),
	.prn(vcc));
defparam \writedata[25] .is_wysiwyg = "true";
defparam \writedata[25] .power_up = "low";

dffeas \writedata[9] (
	.clk(clk_clk),
	.d(writedata_nxt[9]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[9]~q ),
	.prn(vcc));
defparam \writedata[9] .is_wysiwyg = "true";
defparam \writedata[9] .power_up = "low";

dffeas \writedata[18] (
	.clk(clk_clk),
	.d(writedata_nxt[18]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[18]~q ),
	.prn(vcc));
defparam \writedata[18] .is_wysiwyg = "true";
defparam \writedata[18] .power_up = "low";

dffeas \writedata[17] (
	.clk(clk_clk),
	.d(writedata_nxt[17]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[17]~q ),
	.prn(vcc));
defparam \writedata[17] .is_wysiwyg = "true";
defparam \writedata[17] .power_up = "low";

dffeas \readdata[0] (
	.clk(clk_clk),
	.d(\readdata~0_combout ),
	.asdata(\the_processor_cpu_nios2_ocimem|processor_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[0] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_0),
	.prn(vcc));
defparam \readdata[0] .is_wysiwyg = "true";
defparam \readdata[0] .power_up = "low";

dffeas \readdata[16] (
	.clk(clk_clk),
	.d(\the_processor_cpu_nios2_avalon_reg|oci_reg_readdata~0_combout ),
	.asdata(\the_processor_cpu_nios2_ocimem|processor_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[16] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_16),
	.prn(vcc));
defparam \readdata[16] .is_wysiwyg = "true";
defparam \readdata[16] .power_up = "low";

dffeas \readdata[8] (
	.clk(clk_clk),
	.d(\the_processor_cpu_nios2_avalon_reg|oci_reg_readdata~1_combout ),
	.asdata(\the_processor_cpu_nios2_ocimem|processor_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[8] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_8),
	.prn(vcc));
defparam \readdata[8] .is_wysiwyg = "true";
defparam \readdata[8] .power_up = "low";

dffeas \readdata[24] (
	.clk(clk_clk),
	.d(\the_processor_cpu_nios2_avalon_reg|oci_reg_readdata~1_combout ),
	.asdata(\the_processor_cpu_nios2_ocimem|processor_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[24] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_24),
	.prn(vcc));
defparam \readdata[24] .is_wysiwyg = "true";
defparam \readdata[24] .power_up = "low";

dffeas \readdata[5] (
	.clk(clk_clk),
	.d(\the_processor_cpu_nios2_avalon_reg|oci_reg_readdata~1_combout ),
	.asdata(\the_processor_cpu_nios2_ocimem|processor_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[5] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_5),
	.prn(vcc));
defparam \readdata[5] .is_wysiwyg = "true";
defparam \readdata[5] .power_up = "low";

dffeas \readdata[21] (
	.clk(clk_clk),
	.d(\the_processor_cpu_nios2_avalon_reg|oci_reg_readdata~1_combout ),
	.asdata(\the_processor_cpu_nios2_ocimem|processor_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[21] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_21),
	.prn(vcc));
defparam \readdata[21] .is_wysiwyg = "true";
defparam \readdata[21] .power_up = "low";

dffeas \readdata[13] (
	.clk(clk_clk),
	.d(\the_processor_cpu_nios2_avalon_reg|oci_reg_readdata~1_combout ),
	.asdata(\the_processor_cpu_nios2_ocimem|processor_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[13] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_13),
	.prn(vcc));
defparam \readdata[13] .is_wysiwyg = "true";
defparam \readdata[13] .power_up = "low";

dffeas \readdata[29] (
	.clk(clk_clk),
	.d(\the_processor_cpu_nios2_avalon_reg|oci_reg_readdata~1_combout ),
	.asdata(\the_processor_cpu_nios2_ocimem|processor_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[29] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_29),
	.prn(vcc));
defparam \readdata[29] .is_wysiwyg = "true";
defparam \readdata[29] .power_up = "low";

dffeas \readdata[4] (
	.clk(clk_clk),
	.d(\the_processor_cpu_nios2_avalon_reg|oci_reg_readdata~1_combout ),
	.asdata(\the_processor_cpu_nios2_ocimem|processor_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[4] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_4),
	.prn(vcc));
defparam \readdata[4] .is_wysiwyg = "true";
defparam \readdata[4] .power_up = "low";

dffeas \readdata[20] (
	.clk(clk_clk),
	.d(\the_processor_cpu_nios2_avalon_reg|oci_reg_readdata~1_combout ),
	.asdata(\the_processor_cpu_nios2_ocimem|processor_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[20] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_20),
	.prn(vcc));
defparam \readdata[20] .is_wysiwyg = "true";
defparam \readdata[20] .power_up = "low";

dffeas \readdata[12] (
	.clk(clk_clk),
	.d(\the_processor_cpu_nios2_avalon_reg|oci_reg_readdata~1_combout ),
	.asdata(\the_processor_cpu_nios2_ocimem|processor_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[12] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_12),
	.prn(vcc));
defparam \readdata[12] .is_wysiwyg = "true";
defparam \readdata[12] .power_up = "low";

dffeas \readdata[28] (
	.clk(clk_clk),
	.d(\the_processor_cpu_nios2_avalon_reg|oci_reg_readdata~1_combout ),
	.asdata(\the_processor_cpu_nios2_ocimem|processor_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[28] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_28),
	.prn(vcc));
defparam \readdata[28] .is_wysiwyg = "true";
defparam \readdata[28] .power_up = "low";

dffeas \readdata[6] (
	.clk(clk_clk),
	.d(\the_processor_cpu_nios2_avalon_reg|oci_reg_readdata~1_combout ),
	.asdata(\the_processor_cpu_nios2_ocimem|processor_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[6] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_6),
	.prn(vcc));
defparam \readdata[6] .is_wysiwyg = "true";
defparam \readdata[6] .power_up = "low";

dffeas \readdata[22] (
	.clk(clk_clk),
	.d(\the_processor_cpu_nios2_avalon_reg|oci_reg_readdata~1_combout ),
	.asdata(\the_processor_cpu_nios2_ocimem|processor_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[22] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_22),
	.prn(vcc));
defparam \readdata[22] .is_wysiwyg = "true";
defparam \readdata[22] .power_up = "low";

dffeas \readdata[14] (
	.clk(clk_clk),
	.d(\the_processor_cpu_nios2_avalon_reg|oci_reg_readdata~1_combout ),
	.asdata(\the_processor_cpu_nios2_ocimem|processor_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[14] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_14),
	.prn(vcc));
defparam \readdata[14] .is_wysiwyg = "true";
defparam \readdata[14] .power_up = "low";

dffeas \readdata[30] (
	.clk(clk_clk),
	.d(\the_processor_cpu_nios2_avalon_reg|oci_reg_readdata~1_combout ),
	.asdata(\the_processor_cpu_nios2_ocimem|processor_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[30] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_30),
	.prn(vcc));
defparam \readdata[30] .is_wysiwyg = "true";
defparam \readdata[30] .power_up = "low";

dffeas \readdata[7] (
	.clk(clk_clk),
	.d(\the_processor_cpu_nios2_avalon_reg|oci_reg_readdata~1_combout ),
	.asdata(\the_processor_cpu_nios2_ocimem|processor_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[7] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_7),
	.prn(vcc));
defparam \readdata[7] .is_wysiwyg = "true";
defparam \readdata[7] .power_up = "low";

dffeas \readdata[23] (
	.clk(clk_clk),
	.d(\the_processor_cpu_nios2_avalon_reg|oci_reg_readdata~1_combout ),
	.asdata(\the_processor_cpu_nios2_ocimem|processor_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[23] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_23),
	.prn(vcc));
defparam \readdata[23] .is_wysiwyg = "true";
defparam \readdata[23] .power_up = "low";

dffeas \readdata[15] (
	.clk(clk_clk),
	.d(\the_processor_cpu_nios2_avalon_reg|oci_reg_readdata~1_combout ),
	.asdata(\the_processor_cpu_nios2_ocimem|processor_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[15] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_15),
	.prn(vcc));
defparam \readdata[15] .is_wysiwyg = "true";
defparam \readdata[15] .power_up = "low";

dffeas \readdata[31] (
	.clk(clk_clk),
	.d(\the_processor_cpu_nios2_avalon_reg|oci_reg_readdata~1_combout ),
	.asdata(\the_processor_cpu_nios2_ocimem|processor_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[31] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_31),
	.prn(vcc));
defparam \readdata[31] .is_wysiwyg = "true";
defparam \readdata[31] .power_up = "low";

dffeas \readdata[11] (
	.clk(clk_clk),
	.d(\the_processor_cpu_nios2_avalon_reg|oci_reg_readdata~1_combout ),
	.asdata(\the_processor_cpu_nios2_ocimem|processor_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[11] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_11),
	.prn(vcc));
defparam \readdata[11] .is_wysiwyg = "true";
defparam \readdata[11] .power_up = "low";

dffeas \readdata[27] (
	.clk(clk_clk),
	.d(\the_processor_cpu_nios2_avalon_reg|oci_reg_readdata~1_combout ),
	.asdata(\the_processor_cpu_nios2_ocimem|processor_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[27] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_27),
	.prn(vcc));
defparam \readdata[27] .is_wysiwyg = "true";
defparam \readdata[27] .power_up = "low";

dffeas \readdata[10] (
	.clk(clk_clk),
	.d(\the_processor_cpu_nios2_avalon_reg|oci_reg_readdata~1_combout ),
	.asdata(\the_processor_cpu_nios2_ocimem|processor_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[10] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_10),
	.prn(vcc));
defparam \readdata[10] .is_wysiwyg = "true";
defparam \readdata[10] .power_up = "low";

dffeas \readdata[26] (
	.clk(clk_clk),
	.d(\the_processor_cpu_nios2_avalon_reg|oci_reg_readdata~1_combout ),
	.asdata(\the_processor_cpu_nios2_ocimem|processor_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[26] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_26),
	.prn(vcc));
defparam \readdata[26] .is_wysiwyg = "true";
defparam \readdata[26] .power_up = "low";

dffeas \readdata[25] (
	.clk(clk_clk),
	.d(\the_processor_cpu_nios2_avalon_reg|oci_reg_readdata~1_combout ),
	.asdata(\the_processor_cpu_nios2_ocimem|processor_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[25] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_25),
	.prn(vcc));
defparam \readdata[25] .is_wysiwyg = "true";
defparam \readdata[25] .power_up = "low";

dffeas \readdata[9] (
	.clk(clk_clk),
	.d(\the_processor_cpu_nios2_avalon_reg|oci_reg_readdata~1_combout ),
	.asdata(\the_processor_cpu_nios2_ocimem|processor_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[9] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_9),
	.prn(vcc));
defparam \readdata[9] .is_wysiwyg = "true";
defparam \readdata[9] .power_up = "low";

dffeas \readdata[3] (
	.clk(clk_clk),
	.d(\readdata~1_combout ),
	.asdata(\the_processor_cpu_nios2_ocimem|processor_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[3] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_3),
	.prn(vcc));
defparam \readdata[3] .is_wysiwyg = "true";
defparam \readdata[3] .power_up = "low";

dffeas \readdata[19] (
	.clk(clk_clk),
	.d(\the_processor_cpu_nios2_avalon_reg|oci_reg_readdata~1_combout ),
	.asdata(\the_processor_cpu_nios2_ocimem|processor_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[19] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_19),
	.prn(vcc));
defparam \readdata[19] .is_wysiwyg = "true";
defparam \readdata[19] .power_up = "low";

dffeas \readdata[2] (
	.clk(clk_clk),
	.d(\readdata~2_combout ),
	.asdata(\the_processor_cpu_nios2_ocimem|processor_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[2] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_2),
	.prn(vcc));
defparam \readdata[2] .is_wysiwyg = "true";
defparam \readdata[2] .power_up = "low";

dffeas \readdata[18] (
	.clk(clk_clk),
	.d(\the_processor_cpu_nios2_avalon_reg|oci_reg_readdata~1_combout ),
	.asdata(\the_processor_cpu_nios2_ocimem|processor_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[18] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_18),
	.prn(vcc));
defparam \readdata[18] .is_wysiwyg = "true";
defparam \readdata[18] .power_up = "low";

dffeas \readdata[1] (
	.clk(clk_clk),
	.d(\the_processor_cpu_nios2_avalon_reg|oci_reg_readdata[1]~2_combout ),
	.asdata(\the_processor_cpu_nios2_ocimem|processor_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[1] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_1),
	.prn(vcc));
defparam \readdata[1] .is_wysiwyg = "true";
defparam \readdata[1] .power_up = "low";

dffeas \readdata[17] (
	.clk(clk_clk),
	.d(\the_processor_cpu_nios2_avalon_reg|oci_reg_readdata~1_combout ),
	.asdata(\the_processor_cpu_nios2_ocimem|processor_cpu_ociram_sp_ram|the_altsyncram|auto_generated|q_a[17] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_17),
	.prn(vcc));
defparam \readdata[17] .is_wysiwyg = "true";
defparam \readdata[17] .power_up = "low";

cyclonev_lcell_comb \readdata~0 (
	.dataa(!\the_processor_cpu_nios2_avalon_reg|Equal0~1_combout ),
	.datab(!\the_processor_cpu_nios2_oci_debug|monitor_error~q ),
	.datac(!\the_processor_cpu_nios2_avalon_reg|Equal1~0_combout ),
	.datad(!\the_processor_cpu_nios2_avalon_reg|oci_ienable[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\readdata~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata~0 .extended_lut = "off";
defparam \readdata~0 .lut_mask = 64'h27FF27FF27FF27FF;
defparam \readdata~0 .shared_arith = "off";

dffeas \address[8] (
	.clk(clk_clk),
	.d(address_nxt[8]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\address[8]~q ),
	.prn(vcc));
defparam \address[8] .is_wysiwyg = "true";
defparam \address[8] .power_up = "low";

cyclonev_lcell_comb \readdata~1 (
	.dataa(!oci_single_step_mode),
	.datab(!\the_processor_cpu_nios2_avalon_reg|Equal0~1_combout ),
	.datac(!\the_processor_cpu_nios2_avalon_reg|Equal1~0_combout ),
	.datad(!\the_processor_cpu_nios2_avalon_reg|oci_ienable[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\readdata~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata~1 .extended_lut = "off";
defparam \readdata~1 .lut_mask = 64'h47FF47FF47FF47FF;
defparam \readdata~1 .shared_arith = "off";

cyclonev_lcell_comb \readdata~2 (
	.dataa(!\the_processor_cpu_nios2_avalon_reg|Equal0~1_combout ),
	.datab(!\the_processor_cpu_nios2_avalon_reg|Equal1~0_combout ),
	.datac(!\the_processor_cpu_nios2_avalon_reg|oci_ienable[0]~q ),
	.datad(!\the_processor_cpu_nios2_oci_debug|monitor_go~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\readdata~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata~2 .extended_lut = "off";
defparam \readdata~2 .lut_mask = 64'h27FF27FF27FF27FF;
defparam \readdata~2 .shared_arith = "off";

endmodule

module processor_processor_cpu_jtag_debug_module_wrapper (
	break_readreg_0,
	break_readreg_1,
	break_readreg_2,
	MonDReg_2,
	break_readreg_20,
	MonDReg_20,
	break_readreg_19,
	MonDReg_19,
	break_readreg_3,
	break_readreg_16,
	MonDReg_16,
	break_readreg_21,
	MonDReg_21,
	break_readreg_18,
	break_readreg_17,
	MonDReg_17,
	break_readreg_24,
	MonDReg_24,
	break_readreg_4,
	break_readreg_26,
	MonDReg_26,
	break_readreg_25,
	MonDReg_25,
	break_readreg_27,
	MonDReg_27,
	break_readreg_22,
	MonDReg_22,
	MonDReg_13,
	MonDReg_28,
	MonDReg_6,
	MonDReg_14,
	MonDReg_30,
	MonDReg_7,
	MonDReg_23,
	MonDReg_31,
	MonDReg_11,
	MonDReg_10,
	MonDReg_9,
	break_readreg_5,
	break_readreg_28,
	break_readreg_29,
	break_readreg_30,
	break_readreg_31,
	break_readreg_23,
	break_readreg_6,
	break_readreg_15,
	break_readreg_7,
	break_readreg_10,
	break_readreg_14,
	break_readreg_8,
	break_readreg_9,
	break_readreg_13,
	break_readreg_12,
	break_readreg_11,
	sr_0,
	ir_out_0,
	ir_out_1,
	hbreak_enabled,
	MonDReg_0,
	jdo_34,
	jdo_35,
	ir_1,
	ir_0,
	enable_action_strobe,
	take_action_ocimem_a,
	take_action_ocimem_a1,
	take_action_ocimem_a2,
	jdo_21,
	jdo_20,
	monitor_ready,
	MonDReg_1,
	jdo_0,
	jdo_36,
	jdo_37,
	jdo_3,
	jdo_17,
	jdo_19,
	jdo_18,
	jdo_25,
	jdo_1,
	jdo_4,
	jdo_27,
	jdo_26,
	jdo_28,
	monitor_error,
	MonDReg_3,
	jdo_2,
	jdo_5,
	jdo_29,
	jdo_30,
	jdo_31,
	jdo_32,
	jdo_33,
	jdo_23,
	jdo_22,
	MonDReg_18,
	MonDReg_4,
	jdo_6,
	MonDReg_8,
	jdo_16,
	jdo_24,
	MonDReg_5,
	MonDReg_29,
	MonDReg_12,
	MonDReg_15,
	jdo_7,
	resetlatch,
	jdo_11,
	jdo_8,
	jdo_15,
	jdo_9,
	jdo_10,
	jdo_14,
	jdo_13,
	jdo_12,
	altera_internal_jtag,
	altera_internal_jtag1,
	state_4,
	virtual_ir_scan_reg,
	state_3,
	state_8,
	splitter_nodes_receive_1_3,
	irf_reg_0_2,
	irf_reg_1_2,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	break_readreg_0;
input 	break_readreg_1;
input 	break_readreg_2;
input 	MonDReg_2;
input 	break_readreg_20;
input 	MonDReg_20;
input 	break_readreg_19;
input 	MonDReg_19;
input 	break_readreg_3;
input 	break_readreg_16;
input 	MonDReg_16;
input 	break_readreg_21;
input 	MonDReg_21;
input 	break_readreg_18;
input 	break_readreg_17;
input 	MonDReg_17;
input 	break_readreg_24;
input 	MonDReg_24;
input 	break_readreg_4;
input 	break_readreg_26;
input 	MonDReg_26;
input 	break_readreg_25;
input 	MonDReg_25;
input 	break_readreg_27;
input 	MonDReg_27;
input 	break_readreg_22;
input 	MonDReg_22;
input 	MonDReg_13;
input 	MonDReg_28;
input 	MonDReg_6;
input 	MonDReg_14;
input 	MonDReg_30;
input 	MonDReg_7;
input 	MonDReg_23;
input 	MonDReg_31;
input 	MonDReg_11;
input 	MonDReg_10;
input 	MonDReg_9;
input 	break_readreg_5;
input 	break_readreg_28;
input 	break_readreg_29;
input 	break_readreg_30;
input 	break_readreg_31;
input 	break_readreg_23;
input 	break_readreg_6;
input 	break_readreg_15;
input 	break_readreg_7;
input 	break_readreg_10;
input 	break_readreg_14;
input 	break_readreg_8;
input 	break_readreg_9;
input 	break_readreg_13;
input 	break_readreg_12;
input 	break_readreg_11;
output 	sr_0;
output 	ir_out_0;
output 	ir_out_1;
input 	hbreak_enabled;
input 	MonDReg_0;
output 	jdo_34;
output 	jdo_35;
output 	ir_1;
output 	ir_0;
output 	enable_action_strobe;
output 	take_action_ocimem_a;
output 	take_action_ocimem_a1;
output 	take_action_ocimem_a2;
output 	jdo_21;
output 	jdo_20;
input 	monitor_ready;
input 	MonDReg_1;
output 	jdo_0;
output 	jdo_36;
output 	jdo_37;
output 	jdo_3;
output 	jdo_17;
output 	jdo_19;
output 	jdo_18;
output 	jdo_25;
output 	jdo_1;
output 	jdo_4;
output 	jdo_27;
output 	jdo_26;
output 	jdo_28;
input 	monitor_error;
input 	MonDReg_3;
output 	jdo_2;
output 	jdo_5;
output 	jdo_29;
output 	jdo_30;
output 	jdo_31;
output 	jdo_32;
output 	jdo_33;
output 	jdo_23;
output 	jdo_22;
input 	MonDReg_18;
input 	MonDReg_4;
output 	jdo_6;
input 	MonDReg_8;
output 	jdo_16;
output 	jdo_24;
input 	MonDReg_5;
input 	MonDReg_29;
input 	MonDReg_12;
input 	MonDReg_15;
output 	jdo_7;
input 	resetlatch;
output 	jdo_11;
output 	jdo_8;
output 	jdo_15;
output 	jdo_9;
output 	jdo_10;
output 	jdo_14;
output 	jdo_13;
output 	jdo_12;
input 	altera_internal_jtag;
input 	altera_internal_jtag1;
input 	state_4;
input 	virtual_ir_scan_reg;
input 	state_3;
input 	state_8;
input 	splitter_nodes_receive_1_3;
input 	irf_reg_0_2;
input 	irf_reg_1_2;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \the_processor_cpu_jtag_debug_module_tck|sr[1]~q ;
wire \the_processor_cpu_jtag_debug_module_tck|sr[2]~q ;
wire \the_processor_cpu_jtag_debug_module_tck|sr[3]~q ;
wire \the_processor_cpu_jtag_debug_module_tck|sr[21]~q ;
wire \the_processor_cpu_jtag_debug_module_tck|sr[20]~q ;
wire \the_processor_cpu_jtag_debug_module_tck|sr[4]~q ;
wire \the_processor_cpu_jtag_debug_module_tck|sr[17]~q ;
wire \the_processor_cpu_jtag_debug_module_tck|sr[22]~q ;
wire \the_processor_cpu_jtag_debug_module_tck|sr[19]~q ;
wire \the_processor_cpu_jtag_debug_module_tck|sr[18]~q ;
wire \the_processor_cpu_jtag_debug_module_tck|sr[25]~q ;
wire \the_processor_cpu_jtag_debug_module_tck|sr[5]~q ;
wire \the_processor_cpu_jtag_debug_module_tck|sr[27]~q ;
wire \the_processor_cpu_jtag_debug_module_tck|sr[26]~q ;
wire \the_processor_cpu_jtag_debug_module_tck|sr[28]~q ;
wire \the_processor_cpu_jtag_debug_module_tck|sr[23]~q ;
wire \the_processor_cpu_jtag_debug_module_tck|sr[6]~q ;
wire \the_processor_cpu_jtag_debug_module_tck|sr[29]~q ;
wire \the_processor_cpu_jtag_debug_module_tck|sr[30]~q ;
wire \the_processor_cpu_jtag_debug_module_tck|sr[32]~q ;
wire \the_processor_cpu_jtag_debug_module_tck|sr[24]~q ;
wire \the_processor_cpu_jtag_debug_module_tck|sr[16]~q ;
wire \the_processor_cpu_jtag_debug_module_tck|sr[8]~q ;
wire \the_processor_cpu_jtag_debug_module_tck|sr[11]~q ;
wire \the_processor_cpu_jtag_debug_module_tck|sr[9]~q ;
wire \the_processor_cpu_jtag_debug_module_tck|sr[10]~q ;
wire \the_processor_cpu_jtag_debug_module_tck|sr[14]~q ;
wire \the_processor_cpu_jtag_debug_module_tck|sr[13]~q ;
wire \the_processor_cpu_jtag_debug_module_tck|sr[12]~q ;
wire \processor_cpu_jtag_debug_module_phy|virtual_state_sdr~0_combout ;
wire \processor_cpu_jtag_debug_module_phy|virtual_state_uir~combout ;
wire \the_processor_cpu_jtag_debug_module_tck|sr[34]~q ;
wire \the_processor_cpu_jtag_debug_module_tck|sr[35]~q ;
wire \the_processor_cpu_jtag_debug_module_tck|sr[36]~q ;
wire \the_processor_cpu_jtag_debug_module_tck|sr[37]~q ;
wire \processor_cpu_jtag_debug_module_phy|virtual_state_cdr~combout ;
wire \the_processor_cpu_jtag_debug_module_tck|sr[31]~q ;
wire \the_processor_cpu_jtag_debug_module_tck|sr[33]~q ;
wire \processor_cpu_jtag_debug_module_phy|virtual_state_udr~0_combout ;
wire \the_processor_cpu_jtag_debug_module_tck|sr[7]~q ;
wire \the_processor_cpu_jtag_debug_module_tck|sr[15]~q ;


processor_sld_virtual_jtag_basic_1 processor_cpu_jtag_debug_module_phy(
	.virtual_state_sdr(\processor_cpu_jtag_debug_module_phy|virtual_state_sdr~0_combout ),
	.virtual_state_uir1(\processor_cpu_jtag_debug_module_phy|virtual_state_uir~combout ),
	.virtual_state_cdr1(\processor_cpu_jtag_debug_module_phy|virtual_state_cdr~combout ),
	.virtual_state_udr(\processor_cpu_jtag_debug_module_phy|virtual_state_udr~0_combout ),
	.state_4(state_4),
	.virtual_ir_scan_reg(virtual_ir_scan_reg),
	.state_3(state_3),
	.state_8(state_8),
	.splitter_nodes_receive_1_3(splitter_nodes_receive_1_3));

processor_processor_cpu_jtag_debug_module_sysclk the_processor_cpu_jtag_debug_module_sysclk(
	.sr_1(\the_processor_cpu_jtag_debug_module_tck|sr[1]~q ),
	.sr_2(\the_processor_cpu_jtag_debug_module_tck|sr[2]~q ),
	.sr_3(\the_processor_cpu_jtag_debug_module_tck|sr[3]~q ),
	.sr_21(\the_processor_cpu_jtag_debug_module_tck|sr[21]~q ),
	.sr_20(\the_processor_cpu_jtag_debug_module_tck|sr[20]~q ),
	.sr_4(\the_processor_cpu_jtag_debug_module_tck|sr[4]~q ),
	.sr_17(\the_processor_cpu_jtag_debug_module_tck|sr[17]~q ),
	.sr_22(\the_processor_cpu_jtag_debug_module_tck|sr[22]~q ),
	.sr_19(\the_processor_cpu_jtag_debug_module_tck|sr[19]~q ),
	.sr_18(\the_processor_cpu_jtag_debug_module_tck|sr[18]~q ),
	.sr_25(\the_processor_cpu_jtag_debug_module_tck|sr[25]~q ),
	.sr_5(\the_processor_cpu_jtag_debug_module_tck|sr[5]~q ),
	.sr_27(\the_processor_cpu_jtag_debug_module_tck|sr[27]~q ),
	.sr_26(\the_processor_cpu_jtag_debug_module_tck|sr[26]~q ),
	.sr_28(\the_processor_cpu_jtag_debug_module_tck|sr[28]~q ),
	.sr_23(\the_processor_cpu_jtag_debug_module_tck|sr[23]~q ),
	.sr_6(\the_processor_cpu_jtag_debug_module_tck|sr[6]~q ),
	.sr_29(\the_processor_cpu_jtag_debug_module_tck|sr[29]~q ),
	.sr_30(\the_processor_cpu_jtag_debug_module_tck|sr[30]~q ),
	.sr_32(\the_processor_cpu_jtag_debug_module_tck|sr[32]~q ),
	.sr_24(\the_processor_cpu_jtag_debug_module_tck|sr[24]~q ),
	.sr_16(\the_processor_cpu_jtag_debug_module_tck|sr[16]~q ),
	.sr_8(\the_processor_cpu_jtag_debug_module_tck|sr[8]~q ),
	.sr_11(\the_processor_cpu_jtag_debug_module_tck|sr[11]~q ),
	.sr_9(\the_processor_cpu_jtag_debug_module_tck|sr[9]~q ),
	.sr_10(\the_processor_cpu_jtag_debug_module_tck|sr[10]~q ),
	.sr_14(\the_processor_cpu_jtag_debug_module_tck|sr[14]~q ),
	.sr_13(\the_processor_cpu_jtag_debug_module_tck|sr[13]~q ),
	.sr_12(\the_processor_cpu_jtag_debug_module_tck|sr[12]~q ),
	.sr_0(sr_0),
	.virtual_state_uir(\processor_cpu_jtag_debug_module_phy|virtual_state_uir~combout ),
	.jdo_34(jdo_34),
	.jdo_35(jdo_35),
	.ir_1(ir_1),
	.ir_0(ir_0),
	.enable_action_strobe1(enable_action_strobe),
	.take_action_ocimem_a1(take_action_ocimem_a),
	.take_action_ocimem_a2(take_action_ocimem_a1),
	.take_action_ocimem_a3(take_action_ocimem_a2),
	.jdo_21(jdo_21),
	.jdo_20(jdo_20),
	.jdo_0(jdo_0),
	.jdo_36(jdo_36),
	.jdo_37(jdo_37),
	.jdo_3(jdo_3),
	.jdo_17(jdo_17),
	.sr_34(\the_processor_cpu_jtag_debug_module_tck|sr[34]~q ),
	.sr_35(\the_processor_cpu_jtag_debug_module_tck|sr[35]~q ),
	.jdo_19(jdo_19),
	.jdo_18(jdo_18),
	.jdo_25(jdo_25),
	.jdo_1(jdo_1),
	.jdo_4(jdo_4),
	.sr_36(\the_processor_cpu_jtag_debug_module_tck|sr[36]~q ),
	.sr_37(\the_processor_cpu_jtag_debug_module_tck|sr[37]~q ),
	.jdo_27(jdo_27),
	.jdo_26(jdo_26),
	.jdo_28(jdo_28),
	.jdo_2(jdo_2),
	.jdo_5(jdo_5),
	.jdo_29(jdo_29),
	.jdo_30(jdo_30),
	.jdo_31(jdo_31),
	.jdo_32(jdo_32),
	.jdo_33(jdo_33),
	.jdo_23(jdo_23),
	.jdo_22(jdo_22),
	.jdo_6(jdo_6),
	.sr_31(\the_processor_cpu_jtag_debug_module_tck|sr[31]~q ),
	.sr_33(\the_processor_cpu_jtag_debug_module_tck|sr[33]~q ),
	.jdo_16(jdo_16),
	.virtual_state_udr(\processor_cpu_jtag_debug_module_phy|virtual_state_udr~0_combout ),
	.jdo_24(jdo_24),
	.sr_7(\the_processor_cpu_jtag_debug_module_tck|sr[7]~q ),
	.jdo_7(jdo_7),
	.jdo_11(jdo_11),
	.jdo_8(jdo_8),
	.jdo_15(jdo_15),
	.jdo_9(jdo_9),
	.jdo_10(jdo_10),
	.jdo_14(jdo_14),
	.jdo_13(jdo_13),
	.jdo_12(jdo_12),
	.sr_15(\the_processor_cpu_jtag_debug_module_tck|sr[15]~q ),
	.ir_in({irf_reg_1_2,irf_reg_0_2}),
	.clk_clk(clk_clk));

processor_processor_cpu_jtag_debug_module_tck the_processor_cpu_jtag_debug_module_tck(
	.sr_1(\the_processor_cpu_jtag_debug_module_tck|sr[1]~q ),
	.sr_2(\the_processor_cpu_jtag_debug_module_tck|sr[2]~q ),
	.break_readreg_0(break_readreg_0),
	.sr_3(\the_processor_cpu_jtag_debug_module_tck|sr[3]~q ),
	.break_readreg_1(break_readreg_1),
	.sr_21(\the_processor_cpu_jtag_debug_module_tck|sr[21]~q ),
	.sr_20(\the_processor_cpu_jtag_debug_module_tck|sr[20]~q ),
	.sr_4(\the_processor_cpu_jtag_debug_module_tck|sr[4]~q ),
	.break_readreg_2(break_readreg_2),
	.MonDReg_2(MonDReg_2),
	.sr_17(\the_processor_cpu_jtag_debug_module_tck|sr[17]~q ),
	.sr_22(\the_processor_cpu_jtag_debug_module_tck|sr[22]~q ),
	.break_readreg_20(break_readreg_20),
	.MonDReg_20(MonDReg_20),
	.break_readreg_19(break_readreg_19),
	.MonDReg_19(MonDReg_19),
	.sr_19(\the_processor_cpu_jtag_debug_module_tck|sr[19]~q ),
	.sr_18(\the_processor_cpu_jtag_debug_module_tck|sr[18]~q ),
	.sr_25(\the_processor_cpu_jtag_debug_module_tck|sr[25]~q ),
	.sr_5(\the_processor_cpu_jtag_debug_module_tck|sr[5]~q ),
	.break_readreg_3(break_readreg_3),
	.sr_27(\the_processor_cpu_jtag_debug_module_tck|sr[27]~q ),
	.sr_26(\the_processor_cpu_jtag_debug_module_tck|sr[26]~q ),
	.sr_28(\the_processor_cpu_jtag_debug_module_tck|sr[28]~q ),
	.break_readreg_16(break_readreg_16),
	.MonDReg_16(MonDReg_16),
	.sr_23(\the_processor_cpu_jtag_debug_module_tck|sr[23]~q ),
	.break_readreg_21(break_readreg_21),
	.MonDReg_21(MonDReg_21),
	.break_readreg_18(break_readreg_18),
	.break_readreg_17(break_readreg_17),
	.MonDReg_17(MonDReg_17),
	.break_readreg_24(break_readreg_24),
	.MonDReg_24(MonDReg_24),
	.sr_6(\the_processor_cpu_jtag_debug_module_tck|sr[6]~q ),
	.break_readreg_4(break_readreg_4),
	.break_readreg_26(break_readreg_26),
	.MonDReg_26(MonDReg_26),
	.break_readreg_25(break_readreg_25),
	.MonDReg_25(MonDReg_25),
	.sr_29(\the_processor_cpu_jtag_debug_module_tck|sr[29]~q ),
	.break_readreg_27(break_readreg_27),
	.MonDReg_27(MonDReg_27),
	.sr_30(\the_processor_cpu_jtag_debug_module_tck|sr[30]~q ),
	.sr_32(\the_processor_cpu_jtag_debug_module_tck|sr[32]~q ),
	.sr_24(\the_processor_cpu_jtag_debug_module_tck|sr[24]~q ),
	.break_readreg_22(break_readreg_22),
	.MonDReg_22(MonDReg_22),
	.MonDReg_13(MonDReg_13),
	.MonDReg_28(MonDReg_28),
	.MonDReg_6(MonDReg_6),
	.MonDReg_14(MonDReg_14),
	.MonDReg_30(MonDReg_30),
	.MonDReg_7(MonDReg_7),
	.MonDReg_23(MonDReg_23),
	.MonDReg_31(MonDReg_31),
	.MonDReg_11(MonDReg_11),
	.MonDReg_10(MonDReg_10),
	.MonDReg_9(MonDReg_9),
	.break_readreg_5(break_readreg_5),
	.break_readreg_28(break_readreg_28),
	.break_readreg_29(break_readreg_29),
	.break_readreg_30(break_readreg_30),
	.break_readreg_31(break_readreg_31),
	.sr_16(\the_processor_cpu_jtag_debug_module_tck|sr[16]~q ),
	.break_readreg_23(break_readreg_23),
	.sr_8(\the_processor_cpu_jtag_debug_module_tck|sr[8]~q ),
	.break_readreg_6(break_readreg_6),
	.sr_11(\the_processor_cpu_jtag_debug_module_tck|sr[11]~q ),
	.break_readreg_15(break_readreg_15),
	.sr_9(\the_processor_cpu_jtag_debug_module_tck|sr[9]~q ),
	.sr_10(\the_processor_cpu_jtag_debug_module_tck|sr[10]~q ),
	.sr_14(\the_processor_cpu_jtag_debug_module_tck|sr[14]~q ),
	.sr_13(\the_processor_cpu_jtag_debug_module_tck|sr[13]~q ),
	.sr_12(\the_processor_cpu_jtag_debug_module_tck|sr[12]~q ),
	.break_readreg_7(break_readreg_7),
	.break_readreg_10(break_readreg_10),
	.break_readreg_14(break_readreg_14),
	.break_readreg_8(break_readreg_8),
	.break_readreg_9(break_readreg_9),
	.break_readreg_13(break_readreg_13),
	.break_readreg_12(break_readreg_12),
	.break_readreg_11(break_readreg_11),
	.sr_0(sr_0),
	.ir_out_0(ir_out_0),
	.ir_out_1(ir_out_1),
	.virtual_state_sdr(\processor_cpu_jtag_debug_module_phy|virtual_state_sdr~0_combout ),
	.hbreak_enabled(hbreak_enabled),
	.MonDReg_0(MonDReg_0),
	.virtual_state_uir(\processor_cpu_jtag_debug_module_phy|virtual_state_uir~combout ),
	.monitor_ready(monitor_ready),
	.MonDReg_1(MonDReg_1),
	.sr_34(\the_processor_cpu_jtag_debug_module_tck|sr[34]~q ),
	.sr_35(\the_processor_cpu_jtag_debug_module_tck|sr[35]~q ),
	.sr_36(\the_processor_cpu_jtag_debug_module_tck|sr[36]~q ),
	.sr_37(\the_processor_cpu_jtag_debug_module_tck|sr[37]~q ),
	.monitor_error(monitor_error),
	.virtual_state_cdr(\processor_cpu_jtag_debug_module_phy|virtual_state_cdr~combout ),
	.MonDReg_3(MonDReg_3),
	.MonDReg_18(MonDReg_18),
	.MonDReg_4(MonDReg_4),
	.sr_31(\the_processor_cpu_jtag_debug_module_tck|sr[31]~q ),
	.sr_33(\the_processor_cpu_jtag_debug_module_tck|sr[33]~q ),
	.MonDReg_8(MonDReg_8),
	.MonDReg_5(MonDReg_5),
	.MonDReg_29(MonDReg_29),
	.MonDReg_12(MonDReg_12),
	.MonDReg_15(MonDReg_15),
	.sr_7(\the_processor_cpu_jtag_debug_module_tck|sr[7]~q ),
	.resetlatch(resetlatch),
	.sr_15(\the_processor_cpu_jtag_debug_module_tck|sr[15]~q ),
	.altera_internal_jtag(altera_internal_jtag),
	.altera_internal_jtag1(altera_internal_jtag1),
	.state_4(state_4),
	.virtual_ir_scan_reg(virtual_ir_scan_reg),
	.state_3(state_3),
	.splitter_nodes_receive_1_3(splitter_nodes_receive_1_3),
	.irf_reg_0_2(irf_reg_0_2),
	.irf_reg_1_2(irf_reg_1_2));

endmodule

module processor_processor_cpu_jtag_debug_module_sysclk (
	sr_1,
	sr_2,
	sr_3,
	sr_21,
	sr_20,
	sr_4,
	sr_17,
	sr_22,
	sr_19,
	sr_18,
	sr_25,
	sr_5,
	sr_27,
	sr_26,
	sr_28,
	sr_23,
	sr_6,
	sr_29,
	sr_30,
	sr_32,
	sr_24,
	sr_16,
	sr_8,
	sr_11,
	sr_9,
	sr_10,
	sr_14,
	sr_13,
	sr_12,
	sr_0,
	virtual_state_uir,
	jdo_34,
	jdo_35,
	ir_1,
	ir_0,
	enable_action_strobe1,
	take_action_ocimem_a1,
	take_action_ocimem_a2,
	take_action_ocimem_a3,
	jdo_21,
	jdo_20,
	jdo_0,
	jdo_36,
	jdo_37,
	jdo_3,
	jdo_17,
	sr_34,
	sr_35,
	jdo_19,
	jdo_18,
	jdo_25,
	jdo_1,
	jdo_4,
	sr_36,
	sr_37,
	jdo_27,
	jdo_26,
	jdo_28,
	jdo_2,
	jdo_5,
	jdo_29,
	jdo_30,
	jdo_31,
	jdo_32,
	jdo_33,
	jdo_23,
	jdo_22,
	jdo_6,
	sr_31,
	sr_33,
	jdo_16,
	virtual_state_udr,
	jdo_24,
	sr_7,
	jdo_7,
	jdo_11,
	jdo_8,
	jdo_15,
	jdo_9,
	jdo_10,
	jdo_14,
	jdo_13,
	jdo_12,
	sr_15,
	ir_in,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	sr_1;
input 	sr_2;
input 	sr_3;
input 	sr_21;
input 	sr_20;
input 	sr_4;
input 	sr_17;
input 	sr_22;
input 	sr_19;
input 	sr_18;
input 	sr_25;
input 	sr_5;
input 	sr_27;
input 	sr_26;
input 	sr_28;
input 	sr_23;
input 	sr_6;
input 	sr_29;
input 	sr_30;
input 	sr_32;
input 	sr_24;
input 	sr_16;
input 	sr_8;
input 	sr_11;
input 	sr_9;
input 	sr_10;
input 	sr_14;
input 	sr_13;
input 	sr_12;
input 	sr_0;
input 	virtual_state_uir;
output 	jdo_34;
output 	jdo_35;
output 	ir_1;
output 	ir_0;
output 	enable_action_strobe1;
output 	take_action_ocimem_a1;
output 	take_action_ocimem_a2;
output 	take_action_ocimem_a3;
output 	jdo_21;
output 	jdo_20;
output 	jdo_0;
output 	jdo_36;
output 	jdo_37;
output 	jdo_3;
output 	jdo_17;
input 	sr_34;
input 	sr_35;
output 	jdo_19;
output 	jdo_18;
output 	jdo_25;
output 	jdo_1;
output 	jdo_4;
input 	sr_36;
input 	sr_37;
output 	jdo_27;
output 	jdo_26;
output 	jdo_28;
output 	jdo_2;
output 	jdo_5;
output 	jdo_29;
output 	jdo_30;
output 	jdo_31;
output 	jdo_32;
output 	jdo_33;
output 	jdo_23;
output 	jdo_22;
output 	jdo_6;
input 	sr_31;
input 	sr_33;
output 	jdo_16;
input 	virtual_state_udr;
output 	jdo_24;
input 	sr_7;
output 	jdo_7;
output 	jdo_11;
output 	jdo_8;
output 	jdo_15;
output 	jdo_9;
output 	jdo_10;
output 	jdo_14;
output 	jdo_13;
output 	jdo_12;
input 	sr_15;
input 	[1:0] ir_in;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \the_altera_std_synchronizer3|dreg[0]~q ;
wire \the_altera_std_synchronizer4|dreg[0]~q ;
wire \sync2_udr~q ;
wire \update_jdo_strobe~0_combout ;
wire \update_jdo_strobe~q ;
wire \sync2_uir~q ;
wire \jxuir~0_combout ;
wire \jxuir~q ;


processor_altera_std_synchronizer_1 the_altera_std_synchronizer4(
	.din(virtual_state_uir),
	.dreg_0(\the_altera_std_synchronizer4|dreg[0]~q ),
	.clk(clk_clk));

processor_altera_std_synchronizer the_altera_std_synchronizer3(
	.dreg_0(\the_altera_std_synchronizer3|dreg[0]~q ),
	.din(virtual_state_udr),
	.clk(clk_clk));

dffeas \jdo[34] (
	.clk(clk_clk),
	.d(sr_34),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_34),
	.prn(vcc));
defparam \jdo[34] .is_wysiwyg = "true";
defparam \jdo[34] .power_up = "low";

dffeas \jdo[35] (
	.clk(clk_clk),
	.d(sr_35),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_35),
	.prn(vcc));
defparam \jdo[35] .is_wysiwyg = "true";
defparam \jdo[35] .power_up = "low";

dffeas \ir[1] (
	.clk(clk_clk),
	.d(ir_in[1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\jxuir~q ),
	.q(ir_1),
	.prn(vcc));
defparam \ir[1] .is_wysiwyg = "true";
defparam \ir[1] .power_up = "low";

dffeas \ir[0] (
	.clk(clk_clk),
	.d(ir_in[0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\jxuir~q ),
	.q(ir_0),
	.prn(vcc));
defparam \ir[0] .is_wysiwyg = "true";
defparam \ir[0] .power_up = "low";

dffeas enable_action_strobe(
	.clk(clk_clk),
	.d(\update_jdo_strobe~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(enable_action_strobe1),
	.prn(vcc));
defparam enable_action_strobe.is_wysiwyg = "true";
defparam enable_action_strobe.power_up = "low";

cyclonev_lcell_comb \take_action_ocimem_a~0 (
	.dataa(!ir_1),
	.datab(!ir_0),
	.datac(!enable_action_strobe1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(take_action_ocimem_a1),
	.sumout(),
	.cout(),
	.shareout());
defparam \take_action_ocimem_a~0 .extended_lut = "off";
defparam \take_action_ocimem_a~0 .lut_mask = 64'hEFEFEFEFEFEFEFEF;
defparam \take_action_ocimem_a~0 .shared_arith = "off";

cyclonev_lcell_comb \take_action_ocimem_a~1 (
	.dataa(!jdo_35),
	.datab(!take_action_ocimem_a1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(take_action_ocimem_a2),
	.sumout(),
	.cout(),
	.shareout());
defparam \take_action_ocimem_a~1 .extended_lut = "off";
defparam \take_action_ocimem_a~1 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \take_action_ocimem_a~1 .shared_arith = "off";

cyclonev_lcell_comb take_action_ocimem_a(
	.dataa(!jdo_34),
	.datab(!take_action_ocimem_a2),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(take_action_ocimem_a3),
	.sumout(),
	.cout(),
	.shareout());
defparam take_action_ocimem_a.extended_lut = "off";
defparam take_action_ocimem_a.lut_mask = 64'h7777777777777777;
defparam take_action_ocimem_a.shared_arith = "off";

dffeas \jdo[21] (
	.clk(clk_clk),
	.d(sr_21),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_21),
	.prn(vcc));
defparam \jdo[21] .is_wysiwyg = "true";
defparam \jdo[21] .power_up = "low";

dffeas \jdo[20] (
	.clk(clk_clk),
	.d(sr_20),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_20),
	.prn(vcc));
defparam \jdo[20] .is_wysiwyg = "true";
defparam \jdo[20] .power_up = "low";

dffeas \jdo[0] (
	.clk(clk_clk),
	.d(sr_0),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_0),
	.prn(vcc));
defparam \jdo[0] .is_wysiwyg = "true";
defparam \jdo[0] .power_up = "low";

dffeas \jdo[36] (
	.clk(clk_clk),
	.d(sr_36),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_36),
	.prn(vcc));
defparam \jdo[36] .is_wysiwyg = "true";
defparam \jdo[36] .power_up = "low";

dffeas \jdo[37] (
	.clk(clk_clk),
	.d(sr_37),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_37),
	.prn(vcc));
defparam \jdo[37] .is_wysiwyg = "true";
defparam \jdo[37] .power_up = "low";

dffeas \jdo[3] (
	.clk(clk_clk),
	.d(sr_3),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_3),
	.prn(vcc));
defparam \jdo[3] .is_wysiwyg = "true";
defparam \jdo[3] .power_up = "low";

dffeas \jdo[17] (
	.clk(clk_clk),
	.d(sr_17),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_17),
	.prn(vcc));
defparam \jdo[17] .is_wysiwyg = "true";
defparam \jdo[17] .power_up = "low";

dffeas \jdo[19] (
	.clk(clk_clk),
	.d(sr_19),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_19),
	.prn(vcc));
defparam \jdo[19] .is_wysiwyg = "true";
defparam \jdo[19] .power_up = "low";

dffeas \jdo[18] (
	.clk(clk_clk),
	.d(sr_18),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_18),
	.prn(vcc));
defparam \jdo[18] .is_wysiwyg = "true";
defparam \jdo[18] .power_up = "low";

dffeas \jdo[25] (
	.clk(clk_clk),
	.d(sr_25),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_25),
	.prn(vcc));
defparam \jdo[25] .is_wysiwyg = "true";
defparam \jdo[25] .power_up = "low";

dffeas \jdo[1] (
	.clk(clk_clk),
	.d(sr_1),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_1),
	.prn(vcc));
defparam \jdo[1] .is_wysiwyg = "true";
defparam \jdo[1] .power_up = "low";

dffeas \jdo[4] (
	.clk(clk_clk),
	.d(sr_4),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_4),
	.prn(vcc));
defparam \jdo[4] .is_wysiwyg = "true";
defparam \jdo[4] .power_up = "low";

dffeas \jdo[27] (
	.clk(clk_clk),
	.d(sr_27),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_27),
	.prn(vcc));
defparam \jdo[27] .is_wysiwyg = "true";
defparam \jdo[27] .power_up = "low";

dffeas \jdo[26] (
	.clk(clk_clk),
	.d(sr_26),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_26),
	.prn(vcc));
defparam \jdo[26] .is_wysiwyg = "true";
defparam \jdo[26] .power_up = "low";

dffeas \jdo[28] (
	.clk(clk_clk),
	.d(sr_28),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_28),
	.prn(vcc));
defparam \jdo[28] .is_wysiwyg = "true";
defparam \jdo[28] .power_up = "low";

dffeas \jdo[2] (
	.clk(clk_clk),
	.d(sr_2),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_2),
	.prn(vcc));
defparam \jdo[2] .is_wysiwyg = "true";
defparam \jdo[2] .power_up = "low";

dffeas \jdo[5] (
	.clk(clk_clk),
	.d(sr_5),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_5),
	.prn(vcc));
defparam \jdo[5] .is_wysiwyg = "true";
defparam \jdo[5] .power_up = "low";

dffeas \jdo[29] (
	.clk(clk_clk),
	.d(sr_29),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_29),
	.prn(vcc));
defparam \jdo[29] .is_wysiwyg = "true";
defparam \jdo[29] .power_up = "low";

dffeas \jdo[30] (
	.clk(clk_clk),
	.d(sr_30),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_30),
	.prn(vcc));
defparam \jdo[30] .is_wysiwyg = "true";
defparam \jdo[30] .power_up = "low";

dffeas \jdo[31] (
	.clk(clk_clk),
	.d(sr_31),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_31),
	.prn(vcc));
defparam \jdo[31] .is_wysiwyg = "true";
defparam \jdo[31] .power_up = "low";

dffeas \jdo[32] (
	.clk(clk_clk),
	.d(sr_32),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_32),
	.prn(vcc));
defparam \jdo[32] .is_wysiwyg = "true";
defparam \jdo[32] .power_up = "low";

dffeas \jdo[33] (
	.clk(clk_clk),
	.d(sr_33),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_33),
	.prn(vcc));
defparam \jdo[33] .is_wysiwyg = "true";
defparam \jdo[33] .power_up = "low";

dffeas \jdo[23] (
	.clk(clk_clk),
	.d(sr_23),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_23),
	.prn(vcc));
defparam \jdo[23] .is_wysiwyg = "true";
defparam \jdo[23] .power_up = "low";

dffeas \jdo[22] (
	.clk(clk_clk),
	.d(sr_22),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_22),
	.prn(vcc));
defparam \jdo[22] .is_wysiwyg = "true";
defparam \jdo[22] .power_up = "low";

dffeas \jdo[6] (
	.clk(clk_clk),
	.d(sr_6),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_6),
	.prn(vcc));
defparam \jdo[6] .is_wysiwyg = "true";
defparam \jdo[6] .power_up = "low";

dffeas \jdo[16] (
	.clk(clk_clk),
	.d(sr_16),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_16),
	.prn(vcc));
defparam \jdo[16] .is_wysiwyg = "true";
defparam \jdo[16] .power_up = "low";

dffeas \jdo[24] (
	.clk(clk_clk),
	.d(sr_24),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_24),
	.prn(vcc));
defparam \jdo[24] .is_wysiwyg = "true";
defparam \jdo[24] .power_up = "low";

dffeas \jdo[7] (
	.clk(clk_clk),
	.d(sr_7),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_7),
	.prn(vcc));
defparam \jdo[7] .is_wysiwyg = "true";
defparam \jdo[7] .power_up = "low";

dffeas \jdo[11] (
	.clk(clk_clk),
	.d(sr_11),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_11),
	.prn(vcc));
defparam \jdo[11] .is_wysiwyg = "true";
defparam \jdo[11] .power_up = "low";

dffeas \jdo[8] (
	.clk(clk_clk),
	.d(sr_8),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_8),
	.prn(vcc));
defparam \jdo[8] .is_wysiwyg = "true";
defparam \jdo[8] .power_up = "low";

dffeas \jdo[15] (
	.clk(clk_clk),
	.d(sr_15),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_15),
	.prn(vcc));
defparam \jdo[15] .is_wysiwyg = "true";
defparam \jdo[15] .power_up = "low";

dffeas \jdo[9] (
	.clk(clk_clk),
	.d(sr_9),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_9),
	.prn(vcc));
defparam \jdo[9] .is_wysiwyg = "true";
defparam \jdo[9] .power_up = "low";

dffeas \jdo[10] (
	.clk(clk_clk),
	.d(sr_10),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_10),
	.prn(vcc));
defparam \jdo[10] .is_wysiwyg = "true";
defparam \jdo[10] .power_up = "low";

dffeas \jdo[14] (
	.clk(clk_clk),
	.d(sr_14),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_14),
	.prn(vcc));
defparam \jdo[14] .is_wysiwyg = "true";
defparam \jdo[14] .power_up = "low";

dffeas \jdo[13] (
	.clk(clk_clk),
	.d(sr_13),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_13),
	.prn(vcc));
defparam \jdo[13] .is_wysiwyg = "true";
defparam \jdo[13] .power_up = "low";

dffeas \jdo[12] (
	.clk(clk_clk),
	.d(sr_12),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_12),
	.prn(vcc));
defparam \jdo[12] .is_wysiwyg = "true";
defparam \jdo[12] .power_up = "low";

dffeas sync2_udr(
	.clk(clk_clk),
	.d(\the_altera_std_synchronizer3|dreg[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sync2_udr~q ),
	.prn(vcc));
defparam sync2_udr.is_wysiwyg = "true";
defparam sync2_udr.power_up = "low";

cyclonev_lcell_comb \update_jdo_strobe~0 (
	.dataa(!\sync2_udr~q ),
	.datab(!\the_altera_std_synchronizer3|dreg[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\update_jdo_strobe~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \update_jdo_strobe~0 .extended_lut = "off";
defparam \update_jdo_strobe~0 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \update_jdo_strobe~0 .shared_arith = "off";

dffeas update_jdo_strobe(
	.clk(clk_clk),
	.d(\update_jdo_strobe~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\update_jdo_strobe~q ),
	.prn(vcc));
defparam update_jdo_strobe.is_wysiwyg = "true";
defparam update_jdo_strobe.power_up = "low";

dffeas sync2_uir(
	.clk(clk_clk),
	.d(\the_altera_std_synchronizer4|dreg[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sync2_uir~q ),
	.prn(vcc));
defparam sync2_uir.is_wysiwyg = "true";
defparam sync2_uir.power_up = "low";

cyclonev_lcell_comb \jxuir~0 (
	.dataa(!\sync2_uir~q ),
	.datab(!\the_altera_std_synchronizer4|dreg[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\jxuir~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \jxuir~0 .extended_lut = "off";
defparam \jxuir~0 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \jxuir~0 .shared_arith = "off";

dffeas jxuir(
	.clk(clk_clk),
	.d(\jxuir~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\jxuir~q ),
	.prn(vcc));
defparam jxuir.is_wysiwyg = "true";
defparam jxuir.power_up = "low";

endmodule

module processor_altera_std_synchronizer (
	dreg_0,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
output 	dreg_0;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;


dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_0),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

endmodule

module processor_altera_std_synchronizer_1 (
	din,
	dreg_0,
	clk)/* synthesis synthesis_greybox=1 */;
input 	din;
output 	dreg_0;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;


dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_0),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

endmodule

module processor_processor_cpu_jtag_debug_module_tck (
	sr_1,
	sr_2,
	break_readreg_0,
	sr_3,
	break_readreg_1,
	sr_21,
	sr_20,
	sr_4,
	break_readreg_2,
	MonDReg_2,
	sr_17,
	sr_22,
	break_readreg_20,
	MonDReg_20,
	break_readreg_19,
	MonDReg_19,
	sr_19,
	sr_18,
	sr_25,
	sr_5,
	break_readreg_3,
	sr_27,
	sr_26,
	sr_28,
	break_readreg_16,
	MonDReg_16,
	sr_23,
	break_readreg_21,
	MonDReg_21,
	break_readreg_18,
	break_readreg_17,
	MonDReg_17,
	break_readreg_24,
	MonDReg_24,
	sr_6,
	break_readreg_4,
	break_readreg_26,
	MonDReg_26,
	break_readreg_25,
	MonDReg_25,
	sr_29,
	break_readreg_27,
	MonDReg_27,
	sr_30,
	sr_32,
	sr_24,
	break_readreg_22,
	MonDReg_22,
	MonDReg_13,
	MonDReg_28,
	MonDReg_6,
	MonDReg_14,
	MonDReg_30,
	MonDReg_7,
	MonDReg_23,
	MonDReg_31,
	MonDReg_11,
	MonDReg_10,
	MonDReg_9,
	break_readreg_5,
	break_readreg_28,
	break_readreg_29,
	break_readreg_30,
	break_readreg_31,
	sr_16,
	break_readreg_23,
	sr_8,
	break_readreg_6,
	sr_11,
	break_readreg_15,
	sr_9,
	sr_10,
	sr_14,
	sr_13,
	sr_12,
	break_readreg_7,
	break_readreg_10,
	break_readreg_14,
	break_readreg_8,
	break_readreg_9,
	break_readreg_13,
	break_readreg_12,
	break_readreg_11,
	sr_0,
	ir_out_0,
	ir_out_1,
	virtual_state_sdr,
	hbreak_enabled,
	MonDReg_0,
	virtual_state_uir,
	monitor_ready,
	MonDReg_1,
	sr_34,
	sr_35,
	sr_36,
	sr_37,
	monitor_error,
	virtual_state_cdr,
	MonDReg_3,
	MonDReg_18,
	MonDReg_4,
	sr_31,
	sr_33,
	MonDReg_8,
	MonDReg_5,
	MonDReg_29,
	MonDReg_12,
	MonDReg_15,
	sr_7,
	resetlatch,
	sr_15,
	altera_internal_jtag,
	altera_internal_jtag1,
	state_4,
	virtual_ir_scan_reg,
	state_3,
	splitter_nodes_receive_1_3,
	irf_reg_0_2,
	irf_reg_1_2)/* synthesis synthesis_greybox=1 */;
output 	sr_1;
output 	sr_2;
input 	break_readreg_0;
output 	sr_3;
input 	break_readreg_1;
output 	sr_21;
output 	sr_20;
output 	sr_4;
input 	break_readreg_2;
input 	MonDReg_2;
output 	sr_17;
output 	sr_22;
input 	break_readreg_20;
input 	MonDReg_20;
input 	break_readreg_19;
input 	MonDReg_19;
output 	sr_19;
output 	sr_18;
output 	sr_25;
output 	sr_5;
input 	break_readreg_3;
output 	sr_27;
output 	sr_26;
output 	sr_28;
input 	break_readreg_16;
input 	MonDReg_16;
output 	sr_23;
input 	break_readreg_21;
input 	MonDReg_21;
input 	break_readreg_18;
input 	break_readreg_17;
input 	MonDReg_17;
input 	break_readreg_24;
input 	MonDReg_24;
output 	sr_6;
input 	break_readreg_4;
input 	break_readreg_26;
input 	MonDReg_26;
input 	break_readreg_25;
input 	MonDReg_25;
output 	sr_29;
input 	break_readreg_27;
input 	MonDReg_27;
output 	sr_30;
output 	sr_32;
output 	sr_24;
input 	break_readreg_22;
input 	MonDReg_22;
input 	MonDReg_13;
input 	MonDReg_28;
input 	MonDReg_6;
input 	MonDReg_14;
input 	MonDReg_30;
input 	MonDReg_7;
input 	MonDReg_23;
input 	MonDReg_31;
input 	MonDReg_11;
input 	MonDReg_10;
input 	MonDReg_9;
input 	break_readreg_5;
input 	break_readreg_28;
input 	break_readreg_29;
input 	break_readreg_30;
input 	break_readreg_31;
output 	sr_16;
input 	break_readreg_23;
output 	sr_8;
input 	break_readreg_6;
output 	sr_11;
input 	break_readreg_15;
output 	sr_9;
output 	sr_10;
output 	sr_14;
output 	sr_13;
output 	sr_12;
input 	break_readreg_7;
input 	break_readreg_10;
input 	break_readreg_14;
input 	break_readreg_8;
input 	break_readreg_9;
input 	break_readreg_13;
input 	break_readreg_12;
input 	break_readreg_11;
output 	sr_0;
output 	ir_out_0;
output 	ir_out_1;
input 	virtual_state_sdr;
input 	hbreak_enabled;
input 	MonDReg_0;
input 	virtual_state_uir;
input 	monitor_ready;
input 	MonDReg_1;
output 	sr_34;
output 	sr_35;
output 	sr_36;
output 	sr_37;
input 	monitor_error;
input 	virtual_state_cdr;
input 	MonDReg_3;
input 	MonDReg_18;
input 	MonDReg_4;
output 	sr_31;
output 	sr_33;
input 	MonDReg_8;
input 	MonDReg_5;
input 	MonDReg_29;
input 	MonDReg_12;
input 	MonDReg_15;
output 	sr_7;
input 	resetlatch;
output 	sr_15;
input 	altera_internal_jtag;
input 	altera_internal_jtag1;
input 	state_4;
input 	virtual_ir_scan_reg;
input 	state_3;
input 	splitter_nodes_receive_1_3;
input 	irf_reg_0_2;
input 	irf_reg_1_2;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \the_altera_std_synchronizer2|dreg[0]~q ;
wire \the_altera_std_synchronizer1|dreg[0]~q ;
wire \sr~8_combout ;
wire \sr[9]~9_combout ;
wire \sr[9]~10_combout ;
wire \sr~11_combout ;
wire \sr~12_combout ;
wire \sr~16_combout ;
wire \sr[29]~17_combout ;
wire \sr[29]~14_combout ;
wire \sr~18_combout ;
wire \sr~19_combout ;
wire \sr~23_combout ;
wire \sr~24_combout ;
wire \sr~25_combout ;
wire \sr~26_combout ;
wire \sr~27_combout ;
wire \sr~28_combout ;
wire \sr~29_combout ;
wire \sr~30_combout ;
wire \sr~31_combout ;
wire \sr~32_combout ;
wire \sr~33_combout ;
wire \sr~34_combout ;
wire \sr~35_combout ;
wire \sr~40_combout ;
wire \sr~42_combout ;
wire \sr~45_combout ;
wire \sr~46_combout ;
wire \sr~47_combout ;
wire \sr~50_combout ;
wire \sr~51_combout ;
wire \sr~52_combout ;
wire \sr~53_combout ;
wire \sr~54_combout ;
wire \sr~5_combout ;
wire \sr~6_combout ;
wire \DRsize.000~q ;
wire \sr~7_combout ;
wire \Mux37~0_combout ;
wire \sr~13_combout ;
wire \DRsize.100~q ;
wire \sr~56_combout ;
wire \sr~15_combout ;
wire \sr~20_combout ;
wire \sr[36]~21_combout ;
wire \sr~22_combout ;
wire \sr[29]~36_combout ;
wire \sr~37_combout ;
wire \sr~38_combout ;
wire \sr~39_combout ;
wire \sr~41_combout ;
wire \sr~43_combout ;
wire \sr~44_combout ;
wire \sr[29]~55_combout ;
wire \DRsize.010~q ;
wire \sr~48_combout ;
wire \sr~49_combout ;


processor_altera_std_synchronizer_3 the_altera_std_synchronizer2(
	.dreg_0(\the_altera_std_synchronizer2|dreg[0]~q ),
	.din(monitor_ready),
	.clk(altera_internal_jtag));

processor_altera_std_synchronizer_2 the_altera_std_synchronizer1(
	.dreg_0(\the_altera_std_synchronizer1|dreg[0]~q ),
	.din(hbreak_enabled),
	.clk(altera_internal_jtag));

dffeas \sr[1] (
	.clk(altera_internal_jtag),
	.d(\sr~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[9]~9_combout ),
	.sload(gnd),
	.ena(\sr[9]~10_combout ),
	.q(sr_1),
	.prn(vcc));
defparam \sr[1] .is_wysiwyg = "true";
defparam \sr[1] .power_up = "low";

dffeas \sr[2] (
	.clk(altera_internal_jtag),
	.d(\sr~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[9]~9_combout ),
	.sload(gnd),
	.ena(\sr[9]~10_combout ),
	.q(sr_2),
	.prn(vcc));
defparam \sr[2] .is_wysiwyg = "true";
defparam \sr[2] .power_up = "low";

dffeas \sr[3] (
	.clk(altera_internal_jtag),
	.d(\sr~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[9]~9_combout ),
	.sload(gnd),
	.ena(\sr[9]~10_combout ),
	.q(sr_3),
	.prn(vcc));
defparam \sr[3] .is_wysiwyg = "true";
defparam \sr[3] .power_up = "low";

dffeas \sr[21] (
	.clk(altera_internal_jtag),
	.d(\sr~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[29]~17_combout ),
	.sload(gnd),
	.ena(\sr[29]~14_combout ),
	.q(sr_21),
	.prn(vcc));
defparam \sr[21] .is_wysiwyg = "true";
defparam \sr[21] .power_up = "low";

dffeas \sr[20] (
	.clk(altera_internal_jtag),
	.d(\sr~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[29]~17_combout ),
	.sload(gnd),
	.ena(\sr[29]~14_combout ),
	.q(sr_20),
	.prn(vcc));
defparam \sr[20] .is_wysiwyg = "true";
defparam \sr[20] .power_up = "low";

dffeas \sr[4] (
	.clk(altera_internal_jtag),
	.d(\sr~19_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[9]~9_combout ),
	.sload(gnd),
	.ena(\sr[9]~10_combout ),
	.q(sr_4),
	.prn(vcc));
defparam \sr[4] .is_wysiwyg = "true";
defparam \sr[4] .power_up = "low";

dffeas \sr[17] (
	.clk(altera_internal_jtag),
	.d(\sr~23_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[29]~17_combout ),
	.sload(gnd),
	.ena(\sr[29]~14_combout ),
	.q(sr_17),
	.prn(vcc));
defparam \sr[17] .is_wysiwyg = "true";
defparam \sr[17] .power_up = "low";

dffeas \sr[22] (
	.clk(altera_internal_jtag),
	.d(\sr~24_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[29]~17_combout ),
	.sload(gnd),
	.ena(\sr[29]~14_combout ),
	.q(sr_22),
	.prn(vcc));
defparam \sr[22] .is_wysiwyg = "true";
defparam \sr[22] .power_up = "low";

dffeas \sr[19] (
	.clk(altera_internal_jtag),
	.d(\sr~25_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[29]~17_combout ),
	.sload(gnd),
	.ena(\sr[29]~14_combout ),
	.q(sr_19),
	.prn(vcc));
defparam \sr[19] .is_wysiwyg = "true";
defparam \sr[19] .power_up = "low";

dffeas \sr[18] (
	.clk(altera_internal_jtag),
	.d(\sr~26_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[29]~17_combout ),
	.sload(gnd),
	.ena(\sr[29]~14_combout ),
	.q(sr_18),
	.prn(vcc));
defparam \sr[18] .is_wysiwyg = "true";
defparam \sr[18] .power_up = "low";

dffeas \sr[25] (
	.clk(altera_internal_jtag),
	.d(\sr~27_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[29]~17_combout ),
	.sload(gnd),
	.ena(\sr[29]~14_combout ),
	.q(sr_25),
	.prn(vcc));
defparam \sr[25] .is_wysiwyg = "true";
defparam \sr[25] .power_up = "low";

dffeas \sr[5] (
	.clk(altera_internal_jtag),
	.d(\sr~28_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[9]~9_combout ),
	.sload(gnd),
	.ena(\sr[9]~10_combout ),
	.q(sr_5),
	.prn(vcc));
defparam \sr[5] .is_wysiwyg = "true";
defparam \sr[5] .power_up = "low";

dffeas \sr[27] (
	.clk(altera_internal_jtag),
	.d(\sr~29_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[29]~17_combout ),
	.sload(gnd),
	.ena(\sr[29]~14_combout ),
	.q(sr_27),
	.prn(vcc));
defparam \sr[27] .is_wysiwyg = "true";
defparam \sr[27] .power_up = "low";

dffeas \sr[26] (
	.clk(altera_internal_jtag),
	.d(\sr~30_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[29]~17_combout ),
	.sload(gnd),
	.ena(\sr[29]~14_combout ),
	.q(sr_26),
	.prn(vcc));
defparam \sr[26] .is_wysiwyg = "true";
defparam \sr[26] .power_up = "low";

dffeas \sr[28] (
	.clk(altera_internal_jtag),
	.d(\sr~31_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[29]~17_combout ),
	.sload(gnd),
	.ena(\sr[29]~14_combout ),
	.q(sr_28),
	.prn(vcc));
defparam \sr[28] .is_wysiwyg = "true";
defparam \sr[28] .power_up = "low";

dffeas \sr[23] (
	.clk(altera_internal_jtag),
	.d(\sr~32_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[29]~17_combout ),
	.sload(gnd),
	.ena(\sr[29]~14_combout ),
	.q(sr_23),
	.prn(vcc));
defparam \sr[23] .is_wysiwyg = "true";
defparam \sr[23] .power_up = "low";

dffeas \sr[6] (
	.clk(altera_internal_jtag),
	.d(\sr~33_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[9]~9_combout ),
	.sload(gnd),
	.ena(\sr[9]~10_combout ),
	.q(sr_6),
	.prn(vcc));
defparam \sr[6] .is_wysiwyg = "true";
defparam \sr[6] .power_up = "low";

dffeas \sr[29] (
	.clk(altera_internal_jtag),
	.d(\sr~34_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[29]~17_combout ),
	.sload(gnd),
	.ena(\sr[29]~14_combout ),
	.q(sr_29),
	.prn(vcc));
defparam \sr[29] .is_wysiwyg = "true";
defparam \sr[29] .power_up = "low";

dffeas \sr[30] (
	.clk(altera_internal_jtag),
	.d(\sr~35_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[29]~17_combout ),
	.sload(gnd),
	.ena(\sr[29]~14_combout ),
	.q(sr_30),
	.prn(vcc));
defparam \sr[30] .is_wysiwyg = "true";
defparam \sr[30] .power_up = "low";

dffeas \sr[32] (
	.clk(altera_internal_jtag),
	.d(\sr~40_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[29]~17_combout ),
	.sload(gnd),
	.ena(\sr[29]~14_combout ),
	.q(sr_32),
	.prn(vcc));
defparam \sr[32] .is_wysiwyg = "true";
defparam \sr[32] .power_up = "low";

dffeas \sr[24] (
	.clk(altera_internal_jtag),
	.d(\sr~42_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[29]~17_combout ),
	.sload(gnd),
	.ena(\sr[29]~14_combout ),
	.q(sr_24),
	.prn(vcc));
defparam \sr[24] .is_wysiwyg = "true";
defparam \sr[24] .power_up = "low";

dffeas \sr[16] (
	.clk(altera_internal_jtag),
	.d(\sr~45_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[29]~17_combout ),
	.sload(gnd),
	.ena(\sr[29]~14_combout ),
	.q(sr_16),
	.prn(vcc));
defparam \sr[16] .is_wysiwyg = "true";
defparam \sr[16] .power_up = "low";

dffeas \sr[8] (
	.clk(altera_internal_jtag),
	.d(\sr~46_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[9]~9_combout ),
	.sload(gnd),
	.ena(\sr[9]~10_combout ),
	.q(sr_8),
	.prn(vcc));
defparam \sr[8] .is_wysiwyg = "true";
defparam \sr[8] .power_up = "low";

dffeas \sr[11] (
	.clk(altera_internal_jtag),
	.d(\sr~47_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[9]~9_combout ),
	.sload(gnd),
	.ena(\sr[9]~10_combout ),
	.q(sr_11),
	.prn(vcc));
defparam \sr[11] .is_wysiwyg = "true";
defparam \sr[11] .power_up = "low";

dffeas \sr[9] (
	.clk(altera_internal_jtag),
	.d(\sr~50_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[9]~9_combout ),
	.sload(gnd),
	.ena(\sr[9]~10_combout ),
	.q(sr_9),
	.prn(vcc));
defparam \sr[9] .is_wysiwyg = "true";
defparam \sr[9] .power_up = "low";

dffeas \sr[10] (
	.clk(altera_internal_jtag),
	.d(\sr~51_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[9]~9_combout ),
	.sload(gnd),
	.ena(\sr[9]~10_combout ),
	.q(sr_10),
	.prn(vcc));
defparam \sr[10] .is_wysiwyg = "true";
defparam \sr[10] .power_up = "low";

dffeas \sr[14] (
	.clk(altera_internal_jtag),
	.d(\sr~52_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[9]~9_combout ),
	.sload(gnd),
	.ena(\sr[9]~10_combout ),
	.q(sr_14),
	.prn(vcc));
defparam \sr[14] .is_wysiwyg = "true";
defparam \sr[14] .power_up = "low";

dffeas \sr[13] (
	.clk(altera_internal_jtag),
	.d(\sr~53_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[9]~9_combout ),
	.sload(gnd),
	.ena(\sr[9]~10_combout ),
	.q(sr_13),
	.prn(vcc));
defparam \sr[13] .is_wysiwyg = "true";
defparam \sr[13] .power_up = "low";

dffeas \sr[12] (
	.clk(altera_internal_jtag),
	.d(\sr~54_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[9]~9_combout ),
	.sload(gnd),
	.ena(\sr[9]~10_combout ),
	.q(sr_12),
	.prn(vcc));
defparam \sr[12] .is_wysiwyg = "true";
defparam \sr[12] .power_up = "low";

dffeas \sr[0] (
	.clk(altera_internal_jtag),
	.d(\sr~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(sr_0),
	.prn(vcc));
defparam \sr[0] .is_wysiwyg = "true";
defparam \sr[0] .power_up = "low";

dffeas \ir_out[0] (
	.clk(altera_internal_jtag),
	.d(\the_altera_std_synchronizer2|dreg[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(ir_out_0),
	.prn(vcc));
defparam \ir_out[0] .is_wysiwyg = "true";
defparam \ir_out[0] .power_up = "low";

dffeas \ir_out[1] (
	.clk(altera_internal_jtag),
	.d(\the_altera_std_synchronizer1|dreg[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(ir_out_1),
	.prn(vcc));
defparam \ir_out[1] .is_wysiwyg = "true";
defparam \ir_out[1] .power_up = "low";

dffeas \sr[34] (
	.clk(altera_internal_jtag),
	.d(\sr~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[29]~14_combout ),
	.q(sr_34),
	.prn(vcc));
defparam \sr[34] .is_wysiwyg = "true";
defparam \sr[34] .power_up = "low";

dffeas \sr[35] (
	.clk(altera_internal_jtag),
	.d(\sr~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(sr_35),
	.prn(vcc));
defparam \sr[35] .is_wysiwyg = "true";
defparam \sr[35] .power_up = "low";

dffeas \sr[36] (
	.clk(altera_internal_jtag),
	.d(\sr~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[36]~21_combout ),
	.q(sr_36),
	.prn(vcc));
defparam \sr[36] .is_wysiwyg = "true";
defparam \sr[36] .power_up = "low";

dffeas \sr[37] (
	.clk(altera_internal_jtag),
	.d(\sr~22_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[36]~21_combout ),
	.q(sr_37),
	.prn(vcc));
defparam \sr[37] .is_wysiwyg = "true";
defparam \sr[37] .power_up = "low";

dffeas \sr[31] (
	.clk(altera_internal_jtag),
	.d(\sr~39_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(sr_31),
	.prn(vcc));
defparam \sr[31] .is_wysiwyg = "true";
defparam \sr[31] .power_up = "low";

dffeas \sr[33] (
	.clk(altera_internal_jtag),
	.d(\sr~41_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[29]~14_combout ),
	.q(sr_33),
	.prn(vcc));
defparam \sr[33] .is_wysiwyg = "true";
defparam \sr[33] .power_up = "low";

dffeas \sr[7] (
	.clk(altera_internal_jtag),
	.d(\sr~44_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(sr_7),
	.prn(vcc));
defparam \sr[7] .is_wysiwyg = "true";
defparam \sr[7] .power_up = "low";

dffeas \sr[15] (
	.clk(altera_internal_jtag),
	.d(\sr~49_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(sr_15),
	.prn(vcc));
defparam \sr[15] .is_wysiwyg = "true";
defparam \sr[15] .power_up = "low";

cyclonev_lcell_comb \sr~8 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!sr_2),
	.datad(!break_readreg_0),
	.datae(!MonDReg_0),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~8 .extended_lut = "off";
defparam \sr~8 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~8 .shared_arith = "off";

cyclonev_lcell_comb \sr[9]~9 (
	.dataa(!state_4),
	.datab(!virtual_ir_scan_reg),
	.datac(!splitter_nodes_receive_1_3),
	.datad(!irf_reg_0_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr[9]~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr[9]~9 .extended_lut = "off";
defparam \sr[9]~9 .lut_mask = 64'hFBFFFBFFFBFFFBFF;
defparam \sr[9]~9 .shared_arith = "off";

cyclonev_lcell_comb \sr[9]~10 (
	.dataa(!state_4),
	.datab(!virtual_ir_scan_reg),
	.datac(!splitter_nodes_receive_1_3),
	.datad(!state_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr[9]~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr[9]~10 .extended_lut = "off";
defparam \sr[9]~10 .lut_mask = 64'hDFFFDFFFDFFFDFFF;
defparam \sr[9]~10 .shared_arith = "off";

cyclonev_lcell_comb \sr~11 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!sr_3),
	.datad(!break_readreg_1),
	.datae(!MonDReg_1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~11 .extended_lut = "off";
defparam \sr~11 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~11 .shared_arith = "off";

cyclonev_lcell_comb \sr~12 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!sr_4),
	.datad(!break_readreg_2),
	.datae(!MonDReg_2),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~12 .extended_lut = "off";
defparam \sr~12 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~12 .shared_arith = "off";

cyclonev_lcell_comb \sr~16 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!sr_22),
	.datad(!break_readreg_20),
	.datae(!MonDReg_20),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~16 .extended_lut = "off";
defparam \sr~16 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~16 .shared_arith = "off";

cyclonev_lcell_comb \sr[29]~17 (
	.dataa(!state_4),
	.datab(!virtual_ir_scan_reg),
	.datac(!splitter_nodes_receive_1_3),
	.datad(!irf_reg_0_2),
	.datae(!irf_reg_1_2),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr[29]~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr[29]~17 .extended_lut = "off";
defparam \sr[29]~17 .lut_mask = 64'hFFFFFBFFFFFFFBFF;
defparam \sr[29]~17 .shared_arith = "off";

cyclonev_lcell_comb \sr[29]~14 (
	.dataa(!state_4),
	.datab(!virtual_ir_scan_reg),
	.datac(!splitter_nodes_receive_1_3),
	.datad(!state_3),
	.datae(!irf_reg_0_2),
	.dataf(!irf_reg_1_2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr[29]~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr[29]~14 .extended_lut = "off";
defparam \sr[29]~14 .lut_mask = 64'hFFFFFFFFFFFFDFFF;
defparam \sr[29]~14 .shared_arith = "off";

cyclonev_lcell_comb \sr~18 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!sr_21),
	.datad(!break_readreg_19),
	.datae(!MonDReg_19),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~18 .extended_lut = "off";
defparam \sr~18 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~18 .shared_arith = "off";

cyclonev_lcell_comb \sr~19 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!sr_5),
	.datad(!break_readreg_3),
	.datae(!MonDReg_3),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~19 .extended_lut = "off";
defparam \sr~19 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~19 .shared_arith = "off";

cyclonev_lcell_comb \sr~23 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!sr_18),
	.datad(!break_readreg_16),
	.datae(!MonDReg_16),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~23_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~23 .extended_lut = "off";
defparam \sr~23 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~23 .shared_arith = "off";

cyclonev_lcell_comb \sr~24 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!sr_23),
	.datad(!break_readreg_21),
	.datae(!MonDReg_21),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~24_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~24 .extended_lut = "off";
defparam \sr~24 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~24 .shared_arith = "off";

cyclonev_lcell_comb \sr~25 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!sr_20),
	.datad(!break_readreg_18),
	.datae(!MonDReg_18),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~25_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~25 .extended_lut = "off";
defparam \sr~25 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~25 .shared_arith = "off";

cyclonev_lcell_comb \sr~26 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!sr_19),
	.datad(!break_readreg_17),
	.datae(!MonDReg_17),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~26_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~26 .extended_lut = "off";
defparam \sr~26 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~26 .shared_arith = "off";

cyclonev_lcell_comb \sr~27 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!sr_26),
	.datad(!break_readreg_24),
	.datae(!MonDReg_24),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~27_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~27 .extended_lut = "off";
defparam \sr~27 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~27 .shared_arith = "off";

cyclonev_lcell_comb \sr~28 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!sr_6),
	.datad(!break_readreg_4),
	.datae(!MonDReg_4),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~28_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~28 .extended_lut = "off";
defparam \sr~28 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~28 .shared_arith = "off";

cyclonev_lcell_comb \sr~29 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!sr_28),
	.datad(!break_readreg_26),
	.datae(!MonDReg_26),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~29_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~29 .extended_lut = "off";
defparam \sr~29 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~29 .shared_arith = "off";

cyclonev_lcell_comb \sr~30 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!sr_27),
	.datad(!break_readreg_25),
	.datae(!MonDReg_25),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~30_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~30 .extended_lut = "off";
defparam \sr~30 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~30 .shared_arith = "off";

cyclonev_lcell_comb \sr~31 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!sr_29),
	.datad(!break_readreg_27),
	.datae(!MonDReg_27),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~31_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~31 .extended_lut = "off";
defparam \sr~31 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~31 .shared_arith = "off";

cyclonev_lcell_comb \sr~32 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!sr_24),
	.datad(!break_readreg_22),
	.datae(!MonDReg_22),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~32_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~32 .extended_lut = "off";
defparam \sr~32 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~32 .shared_arith = "off";

cyclonev_lcell_comb \sr~33 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!MonDReg_5),
	.datad(!sr_7),
	.datae(!break_readreg_5),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~33_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~33 .extended_lut = "off";
defparam \sr~33 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~33 .shared_arith = "off";

cyclonev_lcell_comb \sr~34 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!sr_30),
	.datad(!MonDReg_28),
	.datae(!break_readreg_28),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~34_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~34 .extended_lut = "off";
defparam \sr~34 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~34 .shared_arith = "off";

cyclonev_lcell_comb \sr~35 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!sr_31),
	.datad(!MonDReg_29),
	.datae(!break_readreg_29),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~35_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~35 .extended_lut = "off";
defparam \sr~35 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~35 .shared_arith = "off";

cyclonev_lcell_comb \sr~40 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!sr_33),
	.datad(!MonDReg_31),
	.datae(!break_readreg_31),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~40_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~40 .extended_lut = "off";
defparam \sr~40 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~40 .shared_arith = "off";

cyclonev_lcell_comb \sr~42 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!sr_25),
	.datad(!MonDReg_23),
	.datae(!break_readreg_23),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~42_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~42 .extended_lut = "off";
defparam \sr~42 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~42 .shared_arith = "off";

cyclonev_lcell_comb \sr~45 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!sr_17),
	.datad(!MonDReg_15),
	.datae(!break_readreg_15),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~45_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~45 .extended_lut = "off";
defparam \sr~45 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~45 .shared_arith = "off";

cyclonev_lcell_comb \sr~46 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!MonDReg_7),
	.datad(!sr_9),
	.datae(!break_readreg_7),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~46_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~46 .extended_lut = "off";
defparam \sr~46 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~46 .shared_arith = "off";

cyclonev_lcell_comb \sr~47 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!MonDReg_10),
	.datad(!sr_12),
	.datae(!break_readreg_10),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~47_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~47 .extended_lut = "off";
defparam \sr~47 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~47 .shared_arith = "off";

cyclonev_lcell_comb \sr~50 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!MonDReg_8),
	.datad(!sr_10),
	.datae(!break_readreg_8),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~50_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~50 .extended_lut = "off";
defparam \sr~50 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~50 .shared_arith = "off";

cyclonev_lcell_comb \sr~51 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!MonDReg_9),
	.datad(!sr_11),
	.datae(!break_readreg_9),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~51_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~51 .extended_lut = "off";
defparam \sr~51 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~51 .shared_arith = "off";

cyclonev_lcell_comb \sr~52 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!MonDReg_13),
	.datad(!sr_15),
	.datae(!break_readreg_13),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~52_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~52 .extended_lut = "off";
defparam \sr~52 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~52 .shared_arith = "off";

cyclonev_lcell_comb \sr~53 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!MonDReg_12),
	.datad(!sr_14),
	.datae(!break_readreg_12),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~53_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~53 .extended_lut = "off";
defparam \sr~53 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~53 .shared_arith = "off";

cyclonev_lcell_comb \sr~54 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_2),
	.datac(!MonDReg_11),
	.datad(!sr_13),
	.datae(!break_readreg_11),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~54_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~54 .extended_lut = "off";
defparam \sr~54 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~54 .shared_arith = "off";

cyclonev_lcell_comb \sr~5 (
	.dataa(!sr_0),
	.datab(!virtual_ir_scan_reg),
	.datac(!splitter_nodes_receive_1_3),
	.datad(!state_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~5 .extended_lut = "off";
defparam \sr~5 .lut_mask = 64'hFFF7FFF7FFF7FFF7;
defparam \sr~5 .shared_arith = "off";

cyclonev_lcell_comb \sr~6 (
	.dataa(!virtual_ir_scan_reg),
	.datab(!splitter_nodes_receive_1_3),
	.datac(!state_3),
	.datad(!\the_altera_std_synchronizer2|dreg[0]~q ),
	.datae(!irf_reg_0_2),
	.dataf(!irf_reg_1_2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~6 .extended_lut = "off";
defparam \sr~6 .lut_mask = 64'hFFFFFFFFFFFFBFFF;
defparam \sr~6 .shared_arith = "off";

dffeas \DRsize.000 (
	.clk(altera_internal_jtag),
	.d(vcc),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(virtual_state_uir),
	.q(\DRsize.000~q ),
	.prn(vcc));
defparam \DRsize.000 .is_wysiwyg = "true";
defparam \DRsize.000 .power_up = "low";

cyclonev_lcell_comb \sr~7 (
	.dataa(!virtual_state_sdr),
	.datab(!\sr~5_combout ),
	.datac(!\sr~6_combout ),
	.datad(!sr_1),
	.datae(!\DRsize.000~q ),
	.dataf(!altera_internal_jtag1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~7 .extended_lut = "off";
defparam \sr~7 .lut_mask = 64'h7FFFBFFFFFFFFFFF;
defparam \sr~7 .shared_arith = "off";

cyclonev_lcell_comb \Mux37~0 (
	.dataa(!irf_reg_0_2),
	.datab(!irf_reg_1_2),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux37~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux37~0 .extended_lut = "off";
defparam \Mux37~0 .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \Mux37~0 .shared_arith = "off";

cyclonev_lcell_comb \sr~13 (
	.dataa(!virtual_state_sdr),
	.datab(!\Mux37~0_combout ),
	.datac(!sr_35),
	.datad(!monitor_error),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~13 .extended_lut = "off";
defparam \sr~13 .lut_mask = 64'h27FF27FF27FF27FF;
defparam \sr~13 .shared_arith = "off";

dffeas \DRsize.100 (
	.clk(altera_internal_jtag),
	.d(\Mux37~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(virtual_state_uir),
	.q(\DRsize.100~q ),
	.prn(vcc));
defparam \DRsize.100 .is_wysiwyg = "true";
defparam \DRsize.100 .power_up = "low";

cyclonev_lcell_comb \sr~56 (
	.dataa(!virtual_state_cdr),
	.datab(!sr_35),
	.datac(!irf_reg_0_2),
	.datad(!irf_reg_1_2),
	.datae(!\the_altera_std_synchronizer1|dreg[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~56_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~56 .extended_lut = "off";
defparam \sr~56 .lut_mask = 64'hB77BFFFFB77BFFFF;
defparam \sr~56 .shared_arith = "off";

cyclonev_lcell_comb \sr~15 (
	.dataa(!virtual_state_sdr),
	.datab(!altera_internal_jtag1),
	.datac(!sr_36),
	.datad(!\DRsize.100~q ),
	.datae(!\sr~56_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~15 .extended_lut = "off";
defparam \sr~15 .lut_mask = 64'h7FBFFFFF7FBFFFFF;
defparam \sr~15 .shared_arith = "off";

cyclonev_lcell_comb \sr~20 (
	.dataa(!state_4),
	.datab(!virtual_ir_scan_reg),
	.datac(!splitter_nodes_receive_1_3),
	.datad(!sr_37),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~20 .extended_lut = "off";
defparam \sr~20 .lut_mask = 64'hDFFFDFFFDFFFDFFF;
defparam \sr~20 .shared_arith = "off";

cyclonev_lcell_comb \sr[36]~21 (
	.dataa(!state_4),
	.datab(!virtual_ir_scan_reg),
	.datac(!splitter_nodes_receive_1_3),
	.datad(!state_3),
	.datae(!irf_reg_0_2),
	.dataf(!irf_reg_1_2),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr[36]~21_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr[36]~21 .extended_lut = "off";
defparam \sr[36]~21 .lut_mask = 64'hDFFFFFFFFFFFDFFF;
defparam \sr[36]~21 .shared_arith = "off";

cyclonev_lcell_comb \sr~22 (
	.dataa(!state_4),
	.datab(!virtual_ir_scan_reg),
	.datac(!splitter_nodes_receive_1_3),
	.datad(!altera_internal_jtag1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~22_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~22 .extended_lut = "off";
defparam \sr~22 .lut_mask = 64'hDFFFDFFFDFFFDFFF;
defparam \sr~22 .shared_arith = "off";

cyclonev_lcell_comb \sr[29]~36 (
	.dataa(!virtual_ir_scan_reg),
	.datab(!splitter_nodes_receive_1_3),
	.datac(!state_3),
	.datad(!irf_reg_0_2),
	.datae(!irf_reg_1_2),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr[29]~36_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr[29]~36 .extended_lut = "off";
defparam \sr[29]~36 .lut_mask = 64'hFFFFFFBFFFFFFFBF;
defparam \sr[29]~36 .shared_arith = "off";

cyclonev_lcell_comb \sr~37 (
	.dataa(!irf_reg_1_2),
	.datab(!MonDReg_30),
	.datac(!break_readreg_30),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~37_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~37 .extended_lut = "off";
defparam \sr~37 .lut_mask = 64'h2727272727272727;
defparam \sr~37 .shared_arith = "off";

cyclonev_lcell_comb \sr~38 (
	.dataa(!virtual_ir_scan_reg),
	.datab(!splitter_nodes_receive_1_3),
	.datac(!state_3),
	.datad(!irf_reg_0_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~38_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~38 .extended_lut = "off";
defparam \sr~38 .lut_mask = 64'hFFBFFFBFFFBFFFBF;
defparam \sr~38 .shared_arith = "off";

cyclonev_lcell_comb \sr~39 (
	.dataa(!virtual_state_sdr),
	.datab(!\sr[29]~36_combout ),
	.datac(!sr_31),
	.datad(!sr_32),
	.datae(!\sr~37_combout ),
	.dataf(!\sr~38_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~39_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~39 .extended_lut = "off";
defparam \sr~39 .lut_mask = 64'h8DFFFFFFFFFFFFFF;
defparam \sr~39 .shared_arith = "off";

cyclonev_lcell_comb \sr~41 (
	.dataa(!virtual_state_sdr),
	.datab(!\Mux37~0_combout ),
	.datac(!sr_34),
	.datad(!resetlatch),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~41_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~41 .extended_lut = "off";
defparam \sr~41 .lut_mask = 64'h27FF27FF27FF27FF;
defparam \sr~41 .shared_arith = "off";

cyclonev_lcell_comb \sr~43 (
	.dataa(!irf_reg_1_2),
	.datab(!MonDReg_6),
	.datac(!break_readreg_6),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~43_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~43 .extended_lut = "off";
defparam \sr~43 .lut_mask = 64'h2727272727272727;
defparam \sr~43 .shared_arith = "off";

cyclonev_lcell_comb \sr~44 (
	.dataa(!virtual_state_sdr),
	.datab(!virtual_state_cdr),
	.datac(!irf_reg_0_2),
	.datad(!sr_7),
	.datae(!sr_8),
	.dataf(!\sr~43_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~44_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~44 .extended_lut = "off";
defparam \sr~44 .lut_mask = 64'hF6FFFFFFFFFFFFFF;
defparam \sr~44 .shared_arith = "off";

cyclonev_lcell_comb \sr[29]~55 (
	.dataa(!irf_reg_0_2),
	.datab(!irf_reg_1_2),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr[29]~55_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr[29]~55 .extended_lut = "off";
defparam \sr[29]~55 .lut_mask = 64'h7777777777777777;
defparam \sr[29]~55 .shared_arith = "off";

dffeas \DRsize.010 (
	.clk(altera_internal_jtag),
	.d(\sr[29]~55_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(virtual_state_uir),
	.q(\DRsize.010~q ),
	.prn(vcc));
defparam \DRsize.010 .is_wysiwyg = "true";
defparam \DRsize.010 .power_up = "low";

cyclonev_lcell_comb \sr~48 (
	.dataa(!virtual_state_cdr),
	.datab(!irf_reg_0_2),
	.datac(!irf_reg_1_2),
	.datad(!MonDReg_14),
	.datae(!sr_15),
	.dataf(!break_readreg_14),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~48_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~48 .extended_lut = "off";
defparam \sr~48 .lut_mask = 64'hDEFFFFFFFFFFFFFF;
defparam \sr~48 .shared_arith = "off";

cyclonev_lcell_comb \sr~49 (
	.dataa(!virtual_state_sdr),
	.datab(!altera_internal_jtag1),
	.datac(!sr_16),
	.datad(!\DRsize.010~q ),
	.datae(!\sr~48_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~49_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~49 .extended_lut = "off";
defparam \sr~49 .lut_mask = 64'h7FBFFFFF7FBFFFFF;
defparam \sr~49 .shared_arith = "off";

endmodule

module processor_altera_std_synchronizer_2 (
	dreg_0,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
output 	dreg_0;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;


dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_0),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

endmodule

module processor_altera_std_synchronizer_3 (
	dreg_0,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
output 	dreg_0;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;


dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_0),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

endmodule

module processor_sld_virtual_jtag_basic_1 (
	virtual_state_sdr,
	virtual_state_uir1,
	virtual_state_cdr1,
	virtual_state_udr,
	state_4,
	virtual_ir_scan_reg,
	state_3,
	state_8,
	splitter_nodes_receive_1_3)/* synthesis synthesis_greybox=1 */;
output 	virtual_state_sdr;
output 	virtual_state_uir1;
output 	virtual_state_cdr1;
output 	virtual_state_udr;
input 	state_4;
input 	virtual_ir_scan_reg;
input 	state_3;
input 	state_8;
input 	splitter_nodes_receive_1_3;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb \virtual_state_sdr~0 (
	.dataa(!state_4),
	.datab(!virtual_ir_scan_reg),
	.datac(!splitter_nodes_receive_1_3),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(virtual_state_sdr),
	.sumout(),
	.cout(),
	.shareout());
defparam \virtual_state_sdr~0 .extended_lut = "off";
defparam \virtual_state_sdr~0 .lut_mask = 64'hDFDFDFDFDFDFDFDF;
defparam \virtual_state_sdr~0 .shared_arith = "off";

cyclonev_lcell_comb virtual_state_uir(
	.dataa(!virtual_ir_scan_reg),
	.datab(!splitter_nodes_receive_1_3),
	.datac(!state_8),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(virtual_state_uir1),
	.sumout(),
	.cout(),
	.shareout());
defparam virtual_state_uir.extended_lut = "off";
defparam virtual_state_uir.lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam virtual_state_uir.shared_arith = "off";

cyclonev_lcell_comb virtual_state_cdr(
	.dataa(!virtual_ir_scan_reg),
	.datab(!splitter_nodes_receive_1_3),
	.datac(!state_3),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(virtual_state_cdr1),
	.sumout(),
	.cout(),
	.shareout());
defparam virtual_state_cdr.extended_lut = "off";
defparam virtual_state_cdr.lut_mask = 64'hBFBFBFBFBFBFBFBF;
defparam virtual_state_cdr.shared_arith = "off";

cyclonev_lcell_comb \virtual_state_udr~0 (
	.dataa(!virtual_ir_scan_reg),
	.datab(!splitter_nodes_receive_1_3),
	.datac(!state_8),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(virtual_state_udr),
	.sumout(),
	.cout(),
	.shareout());
defparam \virtual_state_udr~0 .extended_lut = "off";
defparam \virtual_state_udr~0 .lut_mask = 64'hBFBFBFBFBFBFBFBF;
defparam \virtual_state_udr~0 .shared_arith = "off";

endmodule

module processor_processor_cpu_nios2_avalon_reg (
	r_sync_rst,
	write,
	address_8,
	oci_single_step_mode1,
	monitor_ready,
	writedata_3,
	address_0,
	address_3,
	address_2,
	address_1,
	address_7,
	address_6,
	address_5,
	address_4,
	Equal0,
	debugaccess,
	take_action_ocireg,
	oci_ienable_16,
	oci_ienable_1,
	writedata_16,
	Equal1,
	writedata_1,
	oci_ienable_0,
	oci_reg_readdata,
	oci_reg_readdata1,
	oci_reg_readdata_1,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	r_sync_rst;
input 	write;
input 	address_8;
output 	oci_single_step_mode1;
input 	monitor_ready;
input 	writedata_3;
input 	address_0;
input 	address_3;
input 	address_2;
input 	address_1;
input 	address_7;
input 	address_6;
input 	address_5;
input 	address_4;
output 	Equal0;
input 	debugaccess;
output 	take_action_ocireg;
output 	oci_ienable_16;
output 	oci_ienable_1;
input 	writedata_16;
output 	Equal1;
input 	writedata_1;
output 	oci_ienable_0;
output 	oci_reg_readdata;
output 	oci_reg_readdata1;
output 	oci_reg_readdata_1;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \oci_single_step_mode~0_combout ;
wire \Equal0~0_combout ;
wire \oci_ienable[16]~0_combout ;
wire \take_action_oci_intr_mask_reg~0_combout ;
wire \oci_ienable[1]~1_combout ;


dffeas oci_single_step_mode(
	.clk(clk_clk),
	.d(\oci_single_step_mode~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(oci_single_step_mode1),
	.prn(vcc));
defparam oci_single_step_mode.is_wysiwyg = "true";
defparam oci_single_step_mode.power_up = "low";

cyclonev_lcell_comb \Equal0~1 (
	.dataa(!address_0),
	.datab(!address_3),
	.datac(!address_2),
	.datad(!address_1),
	.datae(!\Equal0~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Equal0),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~1 .extended_lut = "off";
defparam \Equal0~1 .lut_mask = 64'hFFFEFFFFFFFEFFFF;
defparam \Equal0~1 .shared_arith = "off";

cyclonev_lcell_comb \take_action_ocireg~0 (
	.dataa(!write),
	.datab(!Equal0),
	.datac(!debugaccess),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(take_action_ocireg),
	.sumout(),
	.cout(),
	.shareout());
defparam \take_action_ocireg~0 .extended_lut = "off";
defparam \take_action_ocireg~0 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \take_action_ocireg~0 .shared_arith = "off";

dffeas \oci_ienable[16] (
	.clk(clk_clk),
	.d(\oci_ienable[16]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_action_oci_intr_mask_reg~0_combout ),
	.q(oci_ienable_16),
	.prn(vcc));
defparam \oci_ienable[16] .is_wysiwyg = "true";
defparam \oci_ienable[16] .power_up = "low";

dffeas \oci_ienable[1] (
	.clk(clk_clk),
	.d(\oci_ienable[1]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_action_oci_intr_mask_reg~0_combout ),
	.q(oci_ienable_1),
	.prn(vcc));
defparam \oci_ienable[1] .is_wysiwyg = "true";
defparam \oci_ienable[1] .power_up = "low";

cyclonev_lcell_comb \Equal1~0 (
	.dataa(!address_0),
	.datab(!address_3),
	.datac(!address_2),
	.datad(!address_1),
	.datae(!\Equal0~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Equal1),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal1~0 .extended_lut = "off";
defparam \Equal1~0 .lut_mask = 64'hFFFDFFFFFFFDFFFF;
defparam \Equal1~0 .shared_arith = "off";

dffeas \oci_ienable[0] (
	.clk(clk_clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_action_oci_intr_mask_reg~0_combout ),
	.q(oci_ienable_0),
	.prn(vcc));
defparam \oci_ienable[0] .is_wysiwyg = "true";
defparam \oci_ienable[0] .power_up = "low";

cyclonev_lcell_comb \oci_reg_readdata~0 (
	.dataa(!oci_ienable_16),
	.datab(!Equal1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(oci_reg_readdata),
	.sumout(),
	.cout(),
	.shareout());
defparam \oci_reg_readdata~0 .extended_lut = "off";
defparam \oci_reg_readdata~0 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \oci_reg_readdata~0 .shared_arith = "off";

cyclonev_lcell_comb \oci_reg_readdata~1 (
	.dataa(!Equal1),
	.datab(!oci_ienable_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(oci_reg_readdata1),
	.sumout(),
	.cout(),
	.shareout());
defparam \oci_reg_readdata~1 .extended_lut = "off";
defparam \oci_reg_readdata~1 .lut_mask = 64'h7777777777777777;
defparam \oci_reg_readdata~1 .shared_arith = "off";

cyclonev_lcell_comb \oci_reg_readdata[1]~2 (
	.dataa(!monitor_ready),
	.datab(!Equal0),
	.datac(!oci_ienable_1),
	.datad(!Equal1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(oci_reg_readdata_1),
	.sumout(),
	.cout(),
	.shareout());
defparam \oci_reg_readdata[1]~2 .extended_lut = "off";
defparam \oci_reg_readdata[1]~2 .lut_mask = 64'hD1FFD1FFD1FFD1FF;
defparam \oci_reg_readdata[1]~2 .shared_arith = "off";

cyclonev_lcell_comb \oci_single_step_mode~0 (
	.dataa(!oci_single_step_mode1),
	.datab(!writedata_3),
	.datac(!take_action_ocireg),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\oci_single_step_mode~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \oci_single_step_mode~0 .extended_lut = "off";
defparam \oci_single_step_mode~0 .lut_mask = 64'h5353535353535353;
defparam \oci_single_step_mode~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal0~0 (
	.dataa(!address_8),
	.datab(!address_7),
	.datac(!address_6),
	.datad(!address_5),
	.datae(!address_4),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~0 .extended_lut = "off";
defparam \Equal0~0 .lut_mask = 64'hFFFFFFFDFFFFFFFD;
defparam \Equal0~0 .shared_arith = "off";

cyclonev_lcell_comb \oci_ienable[16]~0 (
	.dataa(!writedata_16),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\oci_ienable[16]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \oci_ienable[16]~0 .extended_lut = "off";
defparam \oci_ienable[16]~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \oci_ienable[16]~0 .shared_arith = "off";

cyclonev_lcell_comb \take_action_oci_intr_mask_reg~0 (
	.dataa(!write),
	.datab(!debugaccess),
	.datac(!Equal1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\take_action_oci_intr_mask_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \take_action_oci_intr_mask_reg~0 .extended_lut = "off";
defparam \take_action_oci_intr_mask_reg~0 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \take_action_oci_intr_mask_reg~0 .shared_arith = "off";

cyclonev_lcell_comb \oci_ienable[1]~1 (
	.dataa(!writedata_1),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\oci_ienable[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \oci_ienable[1]~1 .extended_lut = "off";
defparam \oci_ienable[1]~1 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \oci_ienable[1]~1 .shared_arith = "off";

endmodule

module processor_processor_cpu_nios2_oci_break (
	break_readreg_0,
	break_readreg_1,
	break_readreg_2,
	break_readreg_20,
	break_readreg_19,
	break_readreg_3,
	break_readreg_16,
	break_readreg_21,
	break_readreg_18,
	break_readreg_17,
	break_readreg_24,
	break_readreg_4,
	break_readreg_26,
	break_readreg_25,
	break_readreg_27,
	break_readreg_22,
	break_readreg_5,
	break_readreg_28,
	break_readreg_29,
	break_readreg_30,
	break_readreg_31,
	break_readreg_23,
	break_readreg_6,
	break_readreg_15,
	break_readreg_7,
	break_readreg_10,
	break_readreg_14,
	break_readreg_8,
	break_readreg_9,
	break_readreg_13,
	break_readreg_12,
	break_readreg_11,
	ir_1,
	ir_0,
	enable_action_strobe,
	jdo_21,
	jdo_20,
	jdo_0,
	jdo_36,
	jdo_37,
	jdo_3,
	jdo_17,
	jdo_19,
	jdo_18,
	jdo_25,
	jdo_1,
	jdo_4,
	jdo_27,
	jdo_26,
	jdo_28,
	jdo_2,
	jdo_5,
	jdo_29,
	jdo_30,
	jdo_31,
	jdo_23,
	jdo_22,
	jdo_6,
	jdo_16,
	jdo_24,
	jdo_7,
	jdo_11,
	jdo_8,
	jdo_15,
	jdo_9,
	jdo_10,
	jdo_14,
	jdo_13,
	jdo_12,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	break_readreg_0;
output 	break_readreg_1;
output 	break_readreg_2;
output 	break_readreg_20;
output 	break_readreg_19;
output 	break_readreg_3;
output 	break_readreg_16;
output 	break_readreg_21;
output 	break_readreg_18;
output 	break_readreg_17;
output 	break_readreg_24;
output 	break_readreg_4;
output 	break_readreg_26;
output 	break_readreg_25;
output 	break_readreg_27;
output 	break_readreg_22;
output 	break_readreg_5;
output 	break_readreg_28;
output 	break_readreg_29;
output 	break_readreg_30;
output 	break_readreg_31;
output 	break_readreg_23;
output 	break_readreg_6;
output 	break_readreg_15;
output 	break_readreg_7;
output 	break_readreg_10;
output 	break_readreg_14;
output 	break_readreg_8;
output 	break_readreg_9;
output 	break_readreg_13;
output 	break_readreg_12;
output 	break_readreg_11;
input 	ir_1;
input 	ir_0;
input 	enable_action_strobe;
input 	jdo_21;
input 	jdo_20;
input 	jdo_0;
input 	jdo_36;
input 	jdo_37;
input 	jdo_3;
input 	jdo_17;
input 	jdo_19;
input 	jdo_18;
input 	jdo_25;
input 	jdo_1;
input 	jdo_4;
input 	jdo_27;
input 	jdo_26;
input 	jdo_28;
input 	jdo_2;
input 	jdo_5;
input 	jdo_29;
input 	jdo_30;
input 	jdo_31;
input 	jdo_23;
input 	jdo_22;
input 	jdo_6;
input 	jdo_16;
input 	jdo_24;
input 	jdo_7;
input 	jdo_11;
input 	jdo_8;
input 	jdo_15;
input 	jdo_9;
input 	jdo_10;
input 	jdo_14;
input 	jdo_13;
input 	jdo_12;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \break_readreg[27]~0_combout ;
wire \break_readreg[27]~1_combout ;


dffeas \break_readreg[0] (
	.clk(clk_clk),
	.d(jdo_0),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[27]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[27]~0_combout ),
	.q(break_readreg_0),
	.prn(vcc));
defparam \break_readreg[0] .is_wysiwyg = "true";
defparam \break_readreg[0] .power_up = "low";

dffeas \break_readreg[1] (
	.clk(clk_clk),
	.d(jdo_1),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[27]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[27]~0_combout ),
	.q(break_readreg_1),
	.prn(vcc));
defparam \break_readreg[1] .is_wysiwyg = "true";
defparam \break_readreg[1] .power_up = "low";

dffeas \break_readreg[2] (
	.clk(clk_clk),
	.d(jdo_2),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[27]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[27]~0_combout ),
	.q(break_readreg_2),
	.prn(vcc));
defparam \break_readreg[2] .is_wysiwyg = "true";
defparam \break_readreg[2] .power_up = "low";

dffeas \break_readreg[20] (
	.clk(clk_clk),
	.d(jdo_20),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[27]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[27]~0_combout ),
	.q(break_readreg_20),
	.prn(vcc));
defparam \break_readreg[20] .is_wysiwyg = "true";
defparam \break_readreg[20] .power_up = "low";

dffeas \break_readreg[19] (
	.clk(clk_clk),
	.d(jdo_19),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[27]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[27]~0_combout ),
	.q(break_readreg_19),
	.prn(vcc));
defparam \break_readreg[19] .is_wysiwyg = "true";
defparam \break_readreg[19] .power_up = "low";

dffeas \break_readreg[3] (
	.clk(clk_clk),
	.d(jdo_3),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[27]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[27]~0_combout ),
	.q(break_readreg_3),
	.prn(vcc));
defparam \break_readreg[3] .is_wysiwyg = "true";
defparam \break_readreg[3] .power_up = "low";

dffeas \break_readreg[16] (
	.clk(clk_clk),
	.d(jdo_16),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[27]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[27]~0_combout ),
	.q(break_readreg_16),
	.prn(vcc));
defparam \break_readreg[16] .is_wysiwyg = "true";
defparam \break_readreg[16] .power_up = "low";

dffeas \break_readreg[21] (
	.clk(clk_clk),
	.d(jdo_21),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[27]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[27]~0_combout ),
	.q(break_readreg_21),
	.prn(vcc));
defparam \break_readreg[21] .is_wysiwyg = "true";
defparam \break_readreg[21] .power_up = "low";

dffeas \break_readreg[18] (
	.clk(clk_clk),
	.d(jdo_18),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[27]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[27]~0_combout ),
	.q(break_readreg_18),
	.prn(vcc));
defparam \break_readreg[18] .is_wysiwyg = "true";
defparam \break_readreg[18] .power_up = "low";

dffeas \break_readreg[17] (
	.clk(clk_clk),
	.d(jdo_17),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[27]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[27]~0_combout ),
	.q(break_readreg_17),
	.prn(vcc));
defparam \break_readreg[17] .is_wysiwyg = "true";
defparam \break_readreg[17] .power_up = "low";

dffeas \break_readreg[24] (
	.clk(clk_clk),
	.d(jdo_24),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[27]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[27]~0_combout ),
	.q(break_readreg_24),
	.prn(vcc));
defparam \break_readreg[24] .is_wysiwyg = "true";
defparam \break_readreg[24] .power_up = "low";

dffeas \break_readreg[4] (
	.clk(clk_clk),
	.d(jdo_4),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[27]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[27]~0_combout ),
	.q(break_readreg_4),
	.prn(vcc));
defparam \break_readreg[4] .is_wysiwyg = "true";
defparam \break_readreg[4] .power_up = "low";

dffeas \break_readreg[26] (
	.clk(clk_clk),
	.d(jdo_26),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[27]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[27]~0_combout ),
	.q(break_readreg_26),
	.prn(vcc));
defparam \break_readreg[26] .is_wysiwyg = "true";
defparam \break_readreg[26] .power_up = "low";

dffeas \break_readreg[25] (
	.clk(clk_clk),
	.d(jdo_25),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[27]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[27]~0_combout ),
	.q(break_readreg_25),
	.prn(vcc));
defparam \break_readreg[25] .is_wysiwyg = "true";
defparam \break_readreg[25] .power_up = "low";

dffeas \break_readreg[27] (
	.clk(clk_clk),
	.d(jdo_27),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[27]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[27]~0_combout ),
	.q(break_readreg_27),
	.prn(vcc));
defparam \break_readreg[27] .is_wysiwyg = "true";
defparam \break_readreg[27] .power_up = "low";

dffeas \break_readreg[22] (
	.clk(clk_clk),
	.d(jdo_22),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[27]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[27]~0_combout ),
	.q(break_readreg_22),
	.prn(vcc));
defparam \break_readreg[22] .is_wysiwyg = "true";
defparam \break_readreg[22] .power_up = "low";

dffeas \break_readreg[5] (
	.clk(clk_clk),
	.d(jdo_5),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[27]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[27]~0_combout ),
	.q(break_readreg_5),
	.prn(vcc));
defparam \break_readreg[5] .is_wysiwyg = "true";
defparam \break_readreg[5] .power_up = "low";

dffeas \break_readreg[28] (
	.clk(clk_clk),
	.d(jdo_28),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[27]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[27]~0_combout ),
	.q(break_readreg_28),
	.prn(vcc));
defparam \break_readreg[28] .is_wysiwyg = "true";
defparam \break_readreg[28] .power_up = "low";

dffeas \break_readreg[29] (
	.clk(clk_clk),
	.d(jdo_29),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[27]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[27]~0_combout ),
	.q(break_readreg_29),
	.prn(vcc));
defparam \break_readreg[29] .is_wysiwyg = "true";
defparam \break_readreg[29] .power_up = "low";

dffeas \break_readreg[30] (
	.clk(clk_clk),
	.d(jdo_30),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[27]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[27]~0_combout ),
	.q(break_readreg_30),
	.prn(vcc));
defparam \break_readreg[30] .is_wysiwyg = "true";
defparam \break_readreg[30] .power_up = "low";

dffeas \break_readreg[31] (
	.clk(clk_clk),
	.d(jdo_31),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[27]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[27]~0_combout ),
	.q(break_readreg_31),
	.prn(vcc));
defparam \break_readreg[31] .is_wysiwyg = "true";
defparam \break_readreg[31] .power_up = "low";

dffeas \break_readreg[23] (
	.clk(clk_clk),
	.d(jdo_23),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[27]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[27]~0_combout ),
	.q(break_readreg_23),
	.prn(vcc));
defparam \break_readreg[23] .is_wysiwyg = "true";
defparam \break_readreg[23] .power_up = "low";

dffeas \break_readreg[6] (
	.clk(clk_clk),
	.d(jdo_6),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[27]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[27]~0_combout ),
	.q(break_readreg_6),
	.prn(vcc));
defparam \break_readreg[6] .is_wysiwyg = "true";
defparam \break_readreg[6] .power_up = "low";

dffeas \break_readreg[15] (
	.clk(clk_clk),
	.d(jdo_15),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[27]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[27]~0_combout ),
	.q(break_readreg_15),
	.prn(vcc));
defparam \break_readreg[15] .is_wysiwyg = "true";
defparam \break_readreg[15] .power_up = "low";

dffeas \break_readreg[7] (
	.clk(clk_clk),
	.d(jdo_7),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[27]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[27]~0_combout ),
	.q(break_readreg_7),
	.prn(vcc));
defparam \break_readreg[7] .is_wysiwyg = "true";
defparam \break_readreg[7] .power_up = "low";

dffeas \break_readreg[10] (
	.clk(clk_clk),
	.d(jdo_10),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[27]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[27]~0_combout ),
	.q(break_readreg_10),
	.prn(vcc));
defparam \break_readreg[10] .is_wysiwyg = "true";
defparam \break_readreg[10] .power_up = "low";

dffeas \break_readreg[14] (
	.clk(clk_clk),
	.d(jdo_14),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[27]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[27]~0_combout ),
	.q(break_readreg_14),
	.prn(vcc));
defparam \break_readreg[14] .is_wysiwyg = "true";
defparam \break_readreg[14] .power_up = "low";

dffeas \break_readreg[8] (
	.clk(clk_clk),
	.d(jdo_8),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[27]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[27]~0_combout ),
	.q(break_readreg_8),
	.prn(vcc));
defparam \break_readreg[8] .is_wysiwyg = "true";
defparam \break_readreg[8] .power_up = "low";

dffeas \break_readreg[9] (
	.clk(clk_clk),
	.d(jdo_9),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[27]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[27]~0_combout ),
	.q(break_readreg_9),
	.prn(vcc));
defparam \break_readreg[9] .is_wysiwyg = "true";
defparam \break_readreg[9] .power_up = "low";

dffeas \break_readreg[13] (
	.clk(clk_clk),
	.d(jdo_13),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[27]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[27]~0_combout ),
	.q(break_readreg_13),
	.prn(vcc));
defparam \break_readreg[13] .is_wysiwyg = "true";
defparam \break_readreg[13] .power_up = "low";

dffeas \break_readreg[12] (
	.clk(clk_clk),
	.d(jdo_12),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[27]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[27]~0_combout ),
	.q(break_readreg_12),
	.prn(vcc));
defparam \break_readreg[12] .is_wysiwyg = "true";
defparam \break_readreg[12] .power_up = "low";

dffeas \break_readreg[11] (
	.clk(clk_clk),
	.d(jdo_11),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[27]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[27]~0_combout ),
	.q(break_readreg_11),
	.prn(vcc));
defparam \break_readreg[11] .is_wysiwyg = "true";
defparam \break_readreg[11] .power_up = "low";

cyclonev_lcell_comb \break_readreg[27]~0 (
	.dataa(!ir_1),
	.datab(!ir_0),
	.datac(!enable_action_strobe),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\break_readreg[27]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \break_readreg[27]~0 .extended_lut = "off";
defparam \break_readreg[27]~0 .lut_mask = 64'hDFDFDFDFDFDFDFDF;
defparam \break_readreg[27]~0 .shared_arith = "off";

cyclonev_lcell_comb \break_readreg[27]~1 (
	.dataa(!jdo_36),
	.datab(!jdo_37),
	.datac(!\break_readreg[27]~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\break_readreg[27]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \break_readreg[27]~1 .extended_lut = "off";
defparam \break_readreg[27]~1 .lut_mask = 64'hEFEFEFEFEFEFEFEF;
defparam \break_readreg[27]~1 .shared_arith = "off";

endmodule

module processor_processor_cpu_nios2_oci_debug (
	r_sync_rst,
	jtag_break1,
	jdo_34,
	jdo_35,
	take_action_ocimem_a,
	take_action_ocimem_a1,
	jdo_21,
	jdo_20,
	monitor_ready1,
	take_action_ocireg,
	jdo_19,
	jdo_18,
	jdo_25,
	writedata_0,
	monitor_error1,
	writedata_1,
	jdo_23,
	monitor_go1,
	jdo_24,
	resetlatch1,
	state_1,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	r_sync_rst;
output 	jtag_break1;
input 	jdo_34;
input 	jdo_35;
input 	take_action_ocimem_a;
input 	take_action_ocimem_a1;
input 	jdo_21;
input 	jdo_20;
output 	monitor_ready1;
input 	take_action_ocireg;
input 	jdo_19;
input 	jdo_18;
input 	jdo_25;
input 	writedata_0;
output 	monitor_error1;
input 	writedata_1;
input 	jdo_23;
output 	monitor_go1;
input 	jdo_24;
output 	resetlatch1;
input 	state_1;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \the_altera_std_synchronizer|dreg[0]~q ;
wire \break_on_reset~0_combout ;
wire \break_on_reset~q ;
wire \jtag_break~0_combout ;
wire \monitor_ready~0_combout ;
wire \monitor_error~0_combout ;
wire \monitor_go~0_combout ;
wire \resetlatch~0_combout ;


processor_altera_std_synchronizer_4 the_altera_std_synchronizer(
	.din(r_sync_rst),
	.dreg_0(\the_altera_std_synchronizer|dreg[0]~q ),
	.clk(clk_clk));

dffeas jtag_break(
	.clk(clk_clk),
	.d(\jtag_break~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(jtag_break1),
	.prn(vcc));
defparam jtag_break.is_wysiwyg = "true";
defparam jtag_break.power_up = "low";

dffeas monitor_ready(
	.clk(clk_clk),
	.d(\monitor_ready~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(monitor_ready1),
	.prn(vcc));
defparam monitor_ready.is_wysiwyg = "true";
defparam monitor_ready.power_up = "low";

dffeas monitor_error(
	.clk(clk_clk),
	.d(\monitor_error~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(monitor_error1),
	.prn(vcc));
defparam monitor_error.is_wysiwyg = "true";
defparam monitor_error.power_up = "low";

dffeas monitor_go(
	.clk(clk_clk),
	.d(\monitor_go~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(monitor_go1),
	.prn(vcc));
defparam monitor_go.is_wysiwyg = "true";
defparam monitor_go.power_up = "low";

dffeas resetlatch(
	.clk(clk_clk),
	.d(\resetlatch~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(resetlatch1),
	.prn(vcc));
defparam resetlatch.is_wysiwyg = "true";
defparam resetlatch.power_up = "low";

cyclonev_lcell_comb \break_on_reset~0 (
	.dataa(!take_action_ocimem_a1),
	.datab(!\break_on_reset~q ),
	.datac(!jdo_19),
	.datad(!jdo_18),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\break_on_reset~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \break_on_reset~0 .extended_lut = "off";
defparam \break_on_reset~0 .lut_mask = 64'hBF1FBF1FBF1FBF1F;
defparam \break_on_reset~0 .shared_arith = "off";

dffeas break_on_reset(
	.clk(clk_clk),
	.d(\break_on_reset~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\break_on_reset~q ),
	.prn(vcc));
defparam break_on_reset.is_wysiwyg = "true";
defparam break_on_reset.power_up = "low";

cyclonev_lcell_comb \jtag_break~0 (
	.dataa(!jtag_break1),
	.datab(!take_action_ocimem_a1),
	.datac(!jdo_21),
	.datad(!jdo_20),
	.datae(!\break_on_reset~q ),
	.dataf(!\the_altera_std_synchronizer|dreg[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\jtag_break~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \jtag_break~0 .extended_lut = "off";
defparam \jtag_break~0 .lut_mask = 64'hFF7FFFFFFFDFFFFF;
defparam \jtag_break~0 .shared_arith = "off";

cyclonev_lcell_comb \monitor_ready~0 (
	.dataa(!take_action_ocimem_a1),
	.datab(!monitor_ready1),
	.datac(!take_action_ocireg),
	.datad(!jdo_25),
	.datae(!writedata_0),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\monitor_ready~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \monitor_ready~0 .extended_lut = "off";
defparam \monitor_ready~0 .lut_mask = 64'hFFBFFFFFFFBFFFFF;
defparam \monitor_ready~0 .shared_arith = "off";

cyclonev_lcell_comb \monitor_error~0 (
	.dataa(!take_action_ocimem_a1),
	.datab(!take_action_ocireg),
	.datac(!jdo_25),
	.datad(!monitor_error1),
	.datae(!writedata_1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\monitor_error~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \monitor_error~0 .extended_lut = "off";
defparam \monitor_error~0 .lut_mask = 64'hFBFFFFFFFBFFFFFF;
defparam \monitor_error~0 .shared_arith = "off";

cyclonev_lcell_comb \monitor_go~0 (
	.dataa(!jdo_34),
	.datab(!jdo_35),
	.datac(!take_action_ocimem_a),
	.datad(!monitor_go1),
	.datae(!jdo_23),
	.dataf(!state_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\monitor_go~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \monitor_go~0 .extended_lut = "off";
defparam \monitor_go~0 .lut_mask = 64'hFFFFFFFFDFFFFFFF;
defparam \monitor_go~0 .shared_arith = "off";

cyclonev_lcell_comb \resetlatch~0 (
	.dataa(!take_action_ocimem_a1),
	.datab(!\the_altera_std_synchronizer|dreg[0]~q ),
	.datac(!jdo_24),
	.datad(!resetlatch1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\resetlatch~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \resetlatch~0 .extended_lut = "off";
defparam \resetlatch~0 .lut_mask = 64'hFBFFFBFFFBFFFBFF;
defparam \resetlatch~0 .shared_arith = "off";

endmodule

module processor_altera_std_synchronizer_4 (
	din,
	dreg_0,
	clk)/* synthesis synthesis_greybox=1 */;
input 	din;
output 	dreg_0;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;


dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_0),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

endmodule

module processor_processor_cpu_nios2_ocimem (
	q_a_0,
	MonDReg_2,
	q_a_1,
	MonDReg_20,
	MonDReg_19,
	q_a_2,
	q_a_16,
	q_a_8,
	q_a_24,
	MonDReg_16,
	MonDReg_21,
	q_a_20,
	q_a_19,
	MonDReg_17,
	q_a_5,
	q_a_21,
	q_a_13,
	q_a_29,
	q_a_4,
	q_a_12,
	q_a_28,
	q_a_6,
	q_a_22,
	q_a_14,
	q_a_30,
	q_a_7,
	q_a_23,
	q_a_15,
	q_a_31,
	q_a_11,
	q_a_27,
	q_a_10,
	q_a_26,
	q_a_25,
	q_a_9,
	q_a_3,
	q_a_18,
	q_a_17,
	MonDReg_24,
	MonDReg_26,
	MonDReg_25,
	MonDReg_27,
	MonDReg_22,
	MonDReg_13,
	MonDReg_28,
	MonDReg_6,
	MonDReg_14,
	MonDReg_30,
	MonDReg_7,
	MonDReg_23,
	MonDReg_31,
	MonDReg_11,
	MonDReg_10,
	MonDReg_9,
	waitrequest1,
	MonDReg_0,
	write,
	address_8,
	read,
	jdo_34,
	jdo_35,
	take_action_ocimem_a,
	take_no_action_ocimem_a,
	take_action_ocimem_a1,
	jdo_21,
	jdo_20,
	MonDReg_1,
	jdo_3,
	jdo_17,
	writedata_3,
	address_0,
	address_3,
	address_2,
	address_1,
	address_7,
	address_6,
	address_5,
	address_4,
	debugaccess,
	jdo_19,
	jdo_18,
	jdo_25,
	writedata_0,
	jdo_4,
	jdo_27,
	jdo_26,
	jdo_28,
	r_early_rst,
	byteenable_0,
	writedata_16,
	MonDReg_3,
	jdo_5,
	writedata_1,
	jdo_29,
	jdo_30,
	jdo_31,
	jdo_32,
	jdo_33,
	jdo_23,
	jdo_22,
	MonDReg_18,
	MonDReg_4,
	jdo_6,
	writedata_2,
	byteenable_2,
	MonDReg_8,
	writedata_8,
	byteenable_1,
	writedata_24,
	byteenable_3,
	jdo_16,
	jdo_24,
	writedata_20,
	writedata_19,
	MonDReg_5,
	writedata_5,
	writedata_21,
	writedata_13,
	MonDReg_29,
	writedata_29,
	writedata_4,
	MonDReg_12,
	writedata_12,
	writedata_28,
	writedata_6,
	writedata_22,
	writedata_14,
	writedata_30,
	writedata_7,
	writedata_23,
	MonDReg_15,
	writedata_15,
	writedata_31,
	writedata_11,
	writedata_27,
	writedata_10,
	writedata_26,
	writedata_25,
	writedata_9,
	writedata_18,
	writedata_17,
	jdo_7,
	jdo_11,
	jdo_8,
	jdo_15,
	jdo_9,
	jdo_10,
	jdo_14,
	jdo_13,
	jdo_12,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	q_a_0;
output 	MonDReg_2;
output 	q_a_1;
output 	MonDReg_20;
output 	MonDReg_19;
output 	q_a_2;
output 	q_a_16;
output 	q_a_8;
output 	q_a_24;
output 	MonDReg_16;
output 	MonDReg_21;
output 	q_a_20;
output 	q_a_19;
output 	MonDReg_17;
output 	q_a_5;
output 	q_a_21;
output 	q_a_13;
output 	q_a_29;
output 	q_a_4;
output 	q_a_12;
output 	q_a_28;
output 	q_a_6;
output 	q_a_22;
output 	q_a_14;
output 	q_a_30;
output 	q_a_7;
output 	q_a_23;
output 	q_a_15;
output 	q_a_31;
output 	q_a_11;
output 	q_a_27;
output 	q_a_10;
output 	q_a_26;
output 	q_a_25;
output 	q_a_9;
output 	q_a_3;
output 	q_a_18;
output 	q_a_17;
output 	MonDReg_24;
output 	MonDReg_26;
output 	MonDReg_25;
output 	MonDReg_27;
output 	MonDReg_22;
output 	MonDReg_13;
output 	MonDReg_28;
output 	MonDReg_6;
output 	MonDReg_14;
output 	MonDReg_30;
output 	MonDReg_7;
output 	MonDReg_23;
output 	MonDReg_31;
output 	MonDReg_11;
output 	MonDReg_10;
output 	MonDReg_9;
output 	waitrequest1;
output 	MonDReg_0;
input 	write;
input 	address_8;
input 	read;
input 	jdo_34;
input 	jdo_35;
input 	take_action_ocimem_a;
input 	take_no_action_ocimem_a;
input 	take_action_ocimem_a1;
input 	jdo_21;
input 	jdo_20;
output 	MonDReg_1;
input 	jdo_3;
input 	jdo_17;
input 	writedata_3;
input 	address_0;
input 	address_3;
input 	address_2;
input 	address_1;
input 	address_7;
input 	address_6;
input 	address_5;
input 	address_4;
input 	debugaccess;
input 	jdo_19;
input 	jdo_18;
input 	jdo_25;
input 	writedata_0;
input 	jdo_4;
input 	jdo_27;
input 	jdo_26;
input 	jdo_28;
input 	r_early_rst;
input 	byteenable_0;
input 	writedata_16;
output 	MonDReg_3;
input 	jdo_5;
input 	writedata_1;
input 	jdo_29;
input 	jdo_30;
input 	jdo_31;
input 	jdo_32;
input 	jdo_33;
input 	jdo_23;
input 	jdo_22;
output 	MonDReg_18;
output 	MonDReg_4;
input 	jdo_6;
input 	writedata_2;
input 	byteenable_2;
output 	MonDReg_8;
input 	writedata_8;
input 	byteenable_1;
input 	writedata_24;
input 	byteenable_3;
input 	jdo_16;
input 	jdo_24;
input 	writedata_20;
input 	writedata_19;
output 	MonDReg_5;
input 	writedata_5;
input 	writedata_21;
input 	writedata_13;
output 	MonDReg_29;
input 	writedata_29;
input 	writedata_4;
output 	MonDReg_12;
input 	writedata_12;
input 	writedata_28;
input 	writedata_6;
input 	writedata_22;
input 	writedata_14;
input 	writedata_30;
input 	writedata_7;
input 	writedata_23;
output 	MonDReg_15;
input 	writedata_15;
input 	writedata_31;
input 	writedata_11;
input 	writedata_27;
input 	writedata_10;
input 	writedata_26;
input 	writedata_25;
input 	writedata_9;
input 	writedata_18;
input 	writedata_17;
input 	jdo_7;
input 	jdo_11;
input 	jdo_8;
input 	jdo_15;
input 	jdo_9;
input 	jdo_10;
input 	jdo_14;
input 	jdo_13;
input 	jdo_12;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \jtag_ram_wr~q ;
wire \ociram_wr_en~0_combout ;
wire \ociram_reset_req~combout ;
wire \ociram_wr_data[0]~0_combout ;
wire \ociram_addr[0]~0_combout ;
wire \ociram_addr[1]~1_combout ;
wire \ociram_addr[2]~2_combout ;
wire \ociram_addr[3]~3_combout ;
wire \ociram_addr[4]~4_combout ;
wire \ociram_addr[5]~5_combout ;
wire \ociram_addr[6]~6_combout ;
wire \ociram_addr[7]~7_combout ;
wire \ociram_byteenable[0]~0_combout ;
wire \ociram_wr_data[1]~1_combout ;
wire \jtag_ram_wr~0_combout ;
wire \ociram_wr_data[2]~2_combout ;
wire \ociram_wr_data[16]~3_combout ;
wire \ociram_byteenable[2]~1_combout ;
wire \ociram_wr_data[8]~4_combout ;
wire \ociram_byteenable[1]~2_combout ;
wire \ociram_wr_data[24]~5_combout ;
wire \ociram_byteenable[3]~3_combout ;
wire \ociram_wr_data[20]~6_combout ;
wire \ociram_wr_data[19]~7_combout ;
wire \ociram_wr_data[5]~8_combout ;
wire \ociram_wr_data[21]~9_combout ;
wire \ociram_wr_data[13]~10_combout ;
wire \ociram_wr_data[29]~11_combout ;
wire \ociram_wr_data[4]~12_combout ;
wire \ociram_wr_data[12]~13_combout ;
wire \ociram_wr_data[28]~14_combout ;
wire \ociram_wr_data[6]~15_combout ;
wire \ociram_wr_data[22]~16_combout ;
wire \ociram_wr_data[14]~17_combout ;
wire \ociram_wr_data[30]~18_combout ;
wire \ociram_wr_data[7]~19_combout ;
wire \ociram_wr_data[23]~20_combout ;
wire \ociram_wr_data[15]~21_combout ;
wire \ociram_wr_data[31]~22_combout ;
wire \ociram_wr_data[11]~23_combout ;
wire \ociram_wr_data[27]~24_combout ;
wire \ociram_wr_data[10]~25_combout ;
wire \ociram_wr_data[26]~26_combout ;
wire \ociram_wr_data[25]~27_combout ;
wire \ociram_wr_data[9]~28_combout ;
wire \ociram_wr_data[3]~29_combout ;
wire \ociram_wr_data[18]~30_combout ;
wire \ociram_wr_data[17]~31_combout ;
wire \Add0~1_wirecell_combout ;
wire \MonAReg[10]~q ;
wire \Add0~9_sumout ;
wire \MonAReg[2]~q ;
wire \Add0~10 ;
wire \Add0~5_sumout ;
wire \MonAReg[3]~q ;
wire \Add0~6 ;
wire \Add0~13_sumout ;
wire \MonAReg[4]~q ;
wire \Add0~14 ;
wire \Add0~21_sumout ;
wire \MonAReg[5]~q ;
wire \Add0~22 ;
wire \Add0~25_sumout ;
wire \MonAReg[6]~q ;
wire \Add0~26 ;
wire \Add0~29_sumout ;
wire \MonAReg[7]~q ;
wire \Add0~30 ;
wire \Add0~33_sumout ;
wire \MonAReg[8]~q ;
wire \Add0~34 ;
wire \Add0~17_sumout ;
wire \MonAReg[9]~q ;
wire \Add0~18 ;
wire \Add0~1_sumout ;
wire \jtag_ram_rd~0_combout ;
wire \MonDReg[0]~0_combout ;
wire \jtag_ram_rd~q ;
wire \jtag_ram_rd_d1~q ;
wire \MonDReg[0]~1_combout ;
wire \jtag_rd~q ;
wire \jtag_rd_d1~q ;
wire \MonDReg[0]~2_combout ;
wire \jtag_ram_access~0_combout ;
wire \jtag_ram_access~q ;
wire \waitrequest~0_combout ;
wire \avalon_ociram_readdata_ready~0_combout ;
wire \avalon_ociram_readdata_ready~q ;
wire \waitrequest~1_combout ;
wire \MonDReg~15_combout ;
wire \Equal0~0_combout ;
wire \MonDReg~3_combout ;
wire \MonDReg~4_combout ;
wire \MonDReg~12_combout ;
wire \MonDReg~5_combout ;
wire \MonDReg~6_combout ;
wire \MonDReg~7_combout ;
wire \MonDReg~14_combout ;
wire \Equal0~1_combout ;
wire \MonDReg~8_combout ;
wire \MonDReg~9_combout ;
wire \MonDReg~10_combout ;
wire \MonDReg~13_combout ;
wire \MonDReg~11_combout ;


processor_processor_cpu_ociram_sp_ram_module processor_cpu_ociram_sp_ram(
	.q_a_0(q_a_0),
	.q_a_1(q_a_1),
	.q_a_2(q_a_2),
	.q_a_16(q_a_16),
	.q_a_8(q_a_8),
	.q_a_24(q_a_24),
	.q_a_20(q_a_20),
	.q_a_19(q_a_19),
	.q_a_5(q_a_5),
	.q_a_21(q_a_21),
	.q_a_13(q_a_13),
	.q_a_29(q_a_29),
	.q_a_4(q_a_4),
	.q_a_12(q_a_12),
	.q_a_28(q_a_28),
	.q_a_6(q_a_6),
	.q_a_22(q_a_22),
	.q_a_14(q_a_14),
	.q_a_30(q_a_30),
	.q_a_7(q_a_7),
	.q_a_23(q_a_23),
	.q_a_15(q_a_15),
	.q_a_31(q_a_31),
	.q_a_11(q_a_11),
	.q_a_27(q_a_27),
	.q_a_10(q_a_10),
	.q_a_26(q_a_26),
	.q_a_25(q_a_25),
	.q_a_9(q_a_9),
	.q_a_3(q_a_3),
	.q_a_18(q_a_18),
	.q_a_17(q_a_17),
	.ociram_wr_en(\ociram_wr_en~0_combout ),
	.ociram_reset_req(\ociram_reset_req~combout ),
	.ociram_wr_data_0(\ociram_wr_data[0]~0_combout ),
	.ociram_addr_0(\ociram_addr[0]~0_combout ),
	.ociram_addr_1(\ociram_addr[1]~1_combout ),
	.ociram_addr_2(\ociram_addr[2]~2_combout ),
	.ociram_addr_3(\ociram_addr[3]~3_combout ),
	.ociram_addr_4(\ociram_addr[4]~4_combout ),
	.ociram_addr_5(\ociram_addr[5]~5_combout ),
	.ociram_addr_6(\ociram_addr[6]~6_combout ),
	.ociram_addr_7(\ociram_addr[7]~7_combout ),
	.ociram_byteenable_0(\ociram_byteenable[0]~0_combout ),
	.ociram_wr_data_1(\ociram_wr_data[1]~1_combout ),
	.ociram_wr_data_2(\ociram_wr_data[2]~2_combout ),
	.ociram_wr_data_16(\ociram_wr_data[16]~3_combout ),
	.ociram_byteenable_2(\ociram_byteenable[2]~1_combout ),
	.ociram_wr_data_8(\ociram_wr_data[8]~4_combout ),
	.ociram_byteenable_1(\ociram_byteenable[1]~2_combout ),
	.ociram_wr_data_24(\ociram_wr_data[24]~5_combout ),
	.ociram_byteenable_3(\ociram_byteenable[3]~3_combout ),
	.ociram_wr_data_20(\ociram_wr_data[20]~6_combout ),
	.ociram_wr_data_19(\ociram_wr_data[19]~7_combout ),
	.ociram_wr_data_5(\ociram_wr_data[5]~8_combout ),
	.ociram_wr_data_21(\ociram_wr_data[21]~9_combout ),
	.ociram_wr_data_13(\ociram_wr_data[13]~10_combout ),
	.ociram_wr_data_29(\ociram_wr_data[29]~11_combout ),
	.ociram_wr_data_4(\ociram_wr_data[4]~12_combout ),
	.ociram_wr_data_12(\ociram_wr_data[12]~13_combout ),
	.ociram_wr_data_28(\ociram_wr_data[28]~14_combout ),
	.ociram_wr_data_6(\ociram_wr_data[6]~15_combout ),
	.ociram_wr_data_22(\ociram_wr_data[22]~16_combout ),
	.ociram_wr_data_14(\ociram_wr_data[14]~17_combout ),
	.ociram_wr_data_30(\ociram_wr_data[30]~18_combout ),
	.ociram_wr_data_7(\ociram_wr_data[7]~19_combout ),
	.ociram_wr_data_23(\ociram_wr_data[23]~20_combout ),
	.ociram_wr_data_15(\ociram_wr_data[15]~21_combout ),
	.ociram_wr_data_31(\ociram_wr_data[31]~22_combout ),
	.ociram_wr_data_11(\ociram_wr_data[11]~23_combout ),
	.ociram_wr_data_27(\ociram_wr_data[27]~24_combout ),
	.ociram_wr_data_10(\ociram_wr_data[10]~25_combout ),
	.ociram_wr_data_26(\ociram_wr_data[26]~26_combout ),
	.ociram_wr_data_25(\ociram_wr_data[25]~27_combout ),
	.ociram_wr_data_9(\ociram_wr_data[9]~28_combout ),
	.ociram_wr_data_3(\ociram_wr_data[3]~29_combout ),
	.ociram_wr_data_18(\ociram_wr_data[18]~30_combout ),
	.ociram_wr_data_17(\ociram_wr_data[17]~31_combout ),
	.clk_clk(clk_clk));

dffeas jtag_ram_wr(
	.clk(clk_clk),
	.d(\jtag_ram_wr~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!take_no_action_ocimem_a),
	.q(\jtag_ram_wr~q ),
	.prn(vcc));
defparam jtag_ram_wr.is_wysiwyg = "true";
defparam jtag_ram_wr.power_up = "low";

cyclonev_lcell_comb \ociram_wr_en~0 (
	.dataa(!write),
	.datab(!address_8),
	.datac(!\jtag_ram_access~q ),
	.datad(!debugaccess),
	.datae(!\jtag_ram_wr~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_en~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_en~0 .extended_lut = "off";
defparam \ociram_wr_en~0 .lut_mask = 64'hC5FFFFFFC5FFFFFF;
defparam \ociram_wr_en~0 .shared_arith = "off";

cyclonev_lcell_comb ociram_reset_req(
	.dataa(!\jtag_ram_access~q ),
	.datab(!r_early_rst),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_reset_req~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam ociram_reset_req.extended_lut = "off";
defparam ociram_reset_req.lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam ociram_reset_req.shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[0]~0 (
	.dataa(!MonDReg_0),
	.datab(!\jtag_ram_access~q ),
	.datac(!writedata_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[0]~0 .extended_lut = "off";
defparam \ociram_wr_data[0]~0 .lut_mask = 64'h4747474747474747;
defparam \ociram_wr_data[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \ociram_addr[0]~0 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!\MonAReg[2]~q ),
	.datac(!address_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_addr[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_addr[0]~0 .extended_lut = "off";
defparam \ociram_addr[0]~0 .lut_mask = 64'h2727272727272727;
defparam \ociram_addr[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \ociram_addr[1]~1 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!\MonAReg[3]~q ),
	.datac(!address_1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_addr[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_addr[1]~1 .extended_lut = "off";
defparam \ociram_addr[1]~1 .lut_mask = 64'h2727272727272727;
defparam \ociram_addr[1]~1 .shared_arith = "off";

cyclonev_lcell_comb \ociram_addr[2]~2 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!\MonAReg[4]~q ),
	.datac(!address_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_addr[2]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_addr[2]~2 .extended_lut = "off";
defparam \ociram_addr[2]~2 .lut_mask = 64'h2727272727272727;
defparam \ociram_addr[2]~2 .shared_arith = "off";

cyclonev_lcell_comb \ociram_addr[3]~3 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!\MonAReg[5]~q ),
	.datac(!address_3),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_addr[3]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_addr[3]~3 .extended_lut = "off";
defparam \ociram_addr[3]~3 .lut_mask = 64'h2727272727272727;
defparam \ociram_addr[3]~3 .shared_arith = "off";

cyclonev_lcell_comb \ociram_addr[4]~4 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!\MonAReg[6]~q ),
	.datac(!address_4),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_addr[4]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_addr[4]~4 .extended_lut = "off";
defparam \ociram_addr[4]~4 .lut_mask = 64'h2727272727272727;
defparam \ociram_addr[4]~4 .shared_arith = "off";

cyclonev_lcell_comb \ociram_addr[5]~5 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!\MonAReg[7]~q ),
	.datac(!address_5),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_addr[5]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_addr[5]~5 .extended_lut = "off";
defparam \ociram_addr[5]~5 .lut_mask = 64'h2727272727272727;
defparam \ociram_addr[5]~5 .shared_arith = "off";

cyclonev_lcell_comb \ociram_addr[6]~6 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!\MonAReg[8]~q ),
	.datac(!address_6),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_addr[6]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_addr[6]~6 .extended_lut = "off";
defparam \ociram_addr[6]~6 .lut_mask = 64'h2727272727272727;
defparam \ociram_addr[6]~6 .shared_arith = "off";

cyclonev_lcell_comb \ociram_addr[7]~7 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!\MonAReg[9]~q ),
	.datac(!address_7),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_addr[7]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_addr[7]~7 .extended_lut = "off";
defparam \ociram_addr[7]~7 .lut_mask = 64'h2727272727272727;
defparam \ociram_addr[7]~7 .shared_arith = "off";

cyclonev_lcell_comb \ociram_byteenable[0]~0 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!byteenable_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_byteenable[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_byteenable[0]~0 .extended_lut = "off";
defparam \ociram_byteenable[0]~0 .lut_mask = 64'h7777777777777777;
defparam \ociram_byteenable[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[1]~1 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_1),
	.datac(!writedata_1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[1]~1 .extended_lut = "off";
defparam \ociram_wr_data[1]~1 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[1]~1 .shared_arith = "off";

cyclonev_lcell_comb \jtag_ram_wr~0 (
	.dataa(!\MonDReg[0]~0_combout ),
	.datab(!\Add0~1_sumout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\jtag_ram_wr~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \jtag_ram_wr~0 .extended_lut = "off";
defparam \jtag_ram_wr~0 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \jtag_ram_wr~0 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[2]~2 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_2),
	.datac(!writedata_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[2]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[2]~2 .extended_lut = "off";
defparam \ociram_wr_data[2]~2 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[2]~2 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[16]~3 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!writedata_16),
	.datac(!MonDReg_16),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[16]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[16]~3 .extended_lut = "off";
defparam \ociram_wr_data[16]~3 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[16]~3 .shared_arith = "off";

cyclonev_lcell_comb \ociram_byteenable[2]~1 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!byteenable_2),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_byteenable[2]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_byteenable[2]~1 .extended_lut = "off";
defparam \ociram_byteenable[2]~1 .lut_mask = 64'h7777777777777777;
defparam \ociram_byteenable[2]~1 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[8]~4 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_8),
	.datac(!writedata_8),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[8]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[8]~4 .extended_lut = "off";
defparam \ociram_wr_data[8]~4 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[8]~4 .shared_arith = "off";

cyclonev_lcell_comb \ociram_byteenable[1]~2 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!byteenable_1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_byteenable[1]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_byteenable[1]~2 .extended_lut = "off";
defparam \ociram_byteenable[1]~2 .lut_mask = 64'h7777777777777777;
defparam \ociram_byteenable[1]~2 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[24]~5 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_24),
	.datac(!writedata_24),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[24]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[24]~5 .extended_lut = "off";
defparam \ociram_wr_data[24]~5 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[24]~5 .shared_arith = "off";

cyclonev_lcell_comb \ociram_byteenable[3]~3 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!byteenable_3),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_byteenable[3]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_byteenable[3]~3 .extended_lut = "off";
defparam \ociram_byteenable[3]~3 .lut_mask = 64'h7777777777777777;
defparam \ociram_byteenable[3]~3 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[20]~6 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_20),
	.datac(!writedata_20),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[20]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[20]~6 .extended_lut = "off";
defparam \ociram_wr_data[20]~6 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[20]~6 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[19]~7 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_19),
	.datac(!writedata_19),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[19]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[19]~7 .extended_lut = "off";
defparam \ociram_wr_data[19]~7 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[19]~7 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[5]~8 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_5),
	.datac(!writedata_5),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[5]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[5]~8 .extended_lut = "off";
defparam \ociram_wr_data[5]~8 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[5]~8 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[21]~9 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_21),
	.datac(!writedata_21),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[21]~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[21]~9 .extended_lut = "off";
defparam \ociram_wr_data[21]~9 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[21]~9 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[13]~10 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_13),
	.datac(!writedata_13),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[13]~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[13]~10 .extended_lut = "off";
defparam \ociram_wr_data[13]~10 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[13]~10 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[29]~11 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_29),
	.datac(!writedata_29),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[29]~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[29]~11 .extended_lut = "off";
defparam \ociram_wr_data[29]~11 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[29]~11 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[4]~12 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_4),
	.datac(!writedata_4),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[4]~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[4]~12 .extended_lut = "off";
defparam \ociram_wr_data[4]~12 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[4]~12 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[12]~13 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_12),
	.datac(!writedata_12),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[12]~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[12]~13 .extended_lut = "off";
defparam \ociram_wr_data[12]~13 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[12]~13 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[28]~14 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_28),
	.datac(!writedata_28),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[28]~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[28]~14 .extended_lut = "off";
defparam \ociram_wr_data[28]~14 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[28]~14 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[6]~15 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_6),
	.datac(!writedata_6),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[6]~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[6]~15 .extended_lut = "off";
defparam \ociram_wr_data[6]~15 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[6]~15 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[22]~16 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_22),
	.datac(!writedata_22),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[22]~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[22]~16 .extended_lut = "off";
defparam \ociram_wr_data[22]~16 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[22]~16 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[14]~17 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_14),
	.datac(!writedata_14),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[14]~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[14]~17 .extended_lut = "off";
defparam \ociram_wr_data[14]~17 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[14]~17 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[30]~18 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_30),
	.datac(!writedata_30),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[30]~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[30]~18 .extended_lut = "off";
defparam \ociram_wr_data[30]~18 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[30]~18 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[7]~19 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_7),
	.datac(!writedata_7),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[7]~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[7]~19 .extended_lut = "off";
defparam \ociram_wr_data[7]~19 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[7]~19 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[23]~20 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_23),
	.datac(!writedata_23),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[23]~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[23]~20 .extended_lut = "off";
defparam \ociram_wr_data[23]~20 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[23]~20 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[15]~21 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_15),
	.datac(!writedata_15),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[15]~21_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[15]~21 .extended_lut = "off";
defparam \ociram_wr_data[15]~21 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[15]~21 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[31]~22 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_31),
	.datac(!writedata_31),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[31]~22_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[31]~22 .extended_lut = "off";
defparam \ociram_wr_data[31]~22 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[31]~22 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[11]~23 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_11),
	.datac(!writedata_11),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[11]~23_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[11]~23 .extended_lut = "off";
defparam \ociram_wr_data[11]~23 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[11]~23 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[27]~24 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_27),
	.datac(!writedata_27),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[27]~24_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[27]~24 .extended_lut = "off";
defparam \ociram_wr_data[27]~24 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[27]~24 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[10]~25 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_10),
	.datac(!writedata_10),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[10]~25_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[10]~25 .extended_lut = "off";
defparam \ociram_wr_data[10]~25 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[10]~25 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[26]~26 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_26),
	.datac(!writedata_26),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[26]~26_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[26]~26 .extended_lut = "off";
defparam \ociram_wr_data[26]~26 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[26]~26 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[25]~27 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_25),
	.datac(!writedata_25),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[25]~27_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[25]~27 .extended_lut = "off";
defparam \ociram_wr_data[25]~27 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[25]~27 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[9]~28 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_9),
	.datac(!writedata_9),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[9]~28_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[9]~28 .extended_lut = "off";
defparam \ociram_wr_data[9]~28 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[9]~28 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[3]~29 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!writedata_3),
	.datac(!MonDReg_3),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[3]~29_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[3]~29 .extended_lut = "off";
defparam \ociram_wr_data[3]~29 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[3]~29 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[18]~30 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_18),
	.datac(!writedata_18),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[18]~30_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[18]~30 .extended_lut = "off";
defparam \ociram_wr_data[18]~30 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[18]~30 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[17]~31 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_17),
	.datac(!writedata_17),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[17]~31_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[17]~31 .extended_lut = "off";
defparam \ociram_wr_data[17]~31 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[17]~31 .shared_arith = "off";

dffeas \MonDReg[2] (
	.clk(clk_clk),
	.d(jdo_5),
	.asdata(q_a_2),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\MonDReg[0]~1_combout ),
	.sload(\MonDReg[0]~0_combout ),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_2),
	.prn(vcc));
defparam \MonDReg[2] .is_wysiwyg = "true";
defparam \MonDReg[2] .power_up = "low";

dffeas \MonDReg[20] (
	.clk(clk_clk),
	.d(jdo_23),
	.asdata(q_a_20),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\MonDReg[0]~1_combout ),
	.sload(\MonDReg[0]~0_combout ),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_20),
	.prn(vcc));
defparam \MonDReg[20] .is_wysiwyg = "true";
defparam \MonDReg[20] .power_up = "low";

dffeas \MonDReg[19] (
	.clk(clk_clk),
	.d(jdo_22),
	.asdata(q_a_19),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\MonDReg[0]~1_combout ),
	.sload(\MonDReg[0]~0_combout ),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_19),
	.prn(vcc));
defparam \MonDReg[19] .is_wysiwyg = "true";
defparam \MonDReg[19] .power_up = "low";

dffeas \MonDReg[16] (
	.clk(clk_clk),
	.d(jdo_19),
	.asdata(q_a_16),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\MonDReg[0]~1_combout ),
	.sload(\MonDReg[0]~0_combout ),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_16),
	.prn(vcc));
defparam \MonDReg[16] .is_wysiwyg = "true";
defparam \MonDReg[16] .power_up = "low";

dffeas \MonDReg[21] (
	.clk(clk_clk),
	.d(jdo_24),
	.asdata(q_a_21),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\MonDReg[0]~1_combout ),
	.sload(\MonDReg[0]~0_combout ),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_21),
	.prn(vcc));
defparam \MonDReg[21] .is_wysiwyg = "true";
defparam \MonDReg[21] .power_up = "low";

dffeas \MonDReg[17] (
	.clk(clk_clk),
	.d(jdo_20),
	.asdata(q_a_17),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\MonDReg[0]~1_combout ),
	.sload(\MonDReg[0]~0_combout ),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_17),
	.prn(vcc));
defparam \MonDReg[17] .is_wysiwyg = "true";
defparam \MonDReg[17] .power_up = "low";

dffeas \MonDReg[24] (
	.clk(clk_clk),
	.d(jdo_27),
	.asdata(q_a_24),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\MonDReg[0]~1_combout ),
	.sload(\MonDReg[0]~0_combout ),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_24),
	.prn(vcc));
defparam \MonDReg[24] .is_wysiwyg = "true";
defparam \MonDReg[24] .power_up = "low";

dffeas \MonDReg[26] (
	.clk(clk_clk),
	.d(jdo_29),
	.asdata(q_a_26),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\MonDReg[0]~1_combout ),
	.sload(\MonDReg[0]~0_combout ),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_26),
	.prn(vcc));
defparam \MonDReg[26] .is_wysiwyg = "true";
defparam \MonDReg[26] .power_up = "low";

dffeas \MonDReg[25] (
	.clk(clk_clk),
	.d(jdo_28),
	.asdata(q_a_25),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\MonDReg[0]~1_combout ),
	.sload(\MonDReg[0]~0_combout ),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_25),
	.prn(vcc));
defparam \MonDReg[25] .is_wysiwyg = "true";
defparam \MonDReg[25] .power_up = "low";

dffeas \MonDReg[27] (
	.clk(clk_clk),
	.d(jdo_30),
	.asdata(q_a_27),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\MonDReg[0]~1_combout ),
	.sload(\MonDReg[0]~0_combout ),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_27),
	.prn(vcc));
defparam \MonDReg[27] .is_wysiwyg = "true";
defparam \MonDReg[27] .power_up = "low";

dffeas \MonDReg[22] (
	.clk(clk_clk),
	.d(jdo_25),
	.asdata(q_a_22),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\MonDReg[0]~1_combout ),
	.sload(\MonDReg[0]~0_combout ),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_22),
	.prn(vcc));
defparam \MonDReg[22] .is_wysiwyg = "true";
defparam \MonDReg[22] .power_up = "low";

dffeas \MonDReg[13] (
	.clk(clk_clk),
	.d(jdo_16),
	.asdata(q_a_13),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\MonDReg[0]~1_combout ),
	.sload(\MonDReg[0]~0_combout ),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_13),
	.prn(vcc));
defparam \MonDReg[13] .is_wysiwyg = "true";
defparam \MonDReg[13] .power_up = "low";

dffeas \MonDReg[28] (
	.clk(clk_clk),
	.d(jdo_31),
	.asdata(q_a_28),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\MonDReg[0]~1_combout ),
	.sload(\MonDReg[0]~0_combout ),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_28),
	.prn(vcc));
defparam \MonDReg[28] .is_wysiwyg = "true";
defparam \MonDReg[28] .power_up = "low";

dffeas \MonDReg[6] (
	.clk(clk_clk),
	.d(jdo_9),
	.asdata(q_a_6),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\MonDReg[0]~1_combout ),
	.sload(\MonDReg[0]~0_combout ),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_6),
	.prn(vcc));
defparam \MonDReg[6] .is_wysiwyg = "true";
defparam \MonDReg[6] .power_up = "low";

dffeas \MonDReg[14] (
	.clk(clk_clk),
	.d(jdo_17),
	.asdata(q_a_14),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\MonDReg[0]~1_combout ),
	.sload(\MonDReg[0]~0_combout ),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_14),
	.prn(vcc));
defparam \MonDReg[14] .is_wysiwyg = "true";
defparam \MonDReg[14] .power_up = "low";

dffeas \MonDReg[30] (
	.clk(clk_clk),
	.d(jdo_33),
	.asdata(q_a_30),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\MonDReg[0]~1_combout ),
	.sload(\MonDReg[0]~0_combout ),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_30),
	.prn(vcc));
defparam \MonDReg[30] .is_wysiwyg = "true";
defparam \MonDReg[30] .power_up = "low";

dffeas \MonDReg[7] (
	.clk(clk_clk),
	.d(jdo_10),
	.asdata(q_a_7),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\MonDReg[0]~1_combout ),
	.sload(\MonDReg[0]~0_combout ),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_7),
	.prn(vcc));
defparam \MonDReg[7] .is_wysiwyg = "true";
defparam \MonDReg[7] .power_up = "low";

dffeas \MonDReg[23] (
	.clk(clk_clk),
	.d(jdo_26),
	.asdata(q_a_23),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\MonDReg[0]~1_combout ),
	.sload(\MonDReg[0]~0_combout ),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_23),
	.prn(vcc));
defparam \MonDReg[23] .is_wysiwyg = "true";
defparam \MonDReg[23] .power_up = "low";

dffeas \MonDReg[31] (
	.clk(clk_clk),
	.d(jdo_34),
	.asdata(q_a_31),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\MonDReg[0]~1_combout ),
	.sload(\MonDReg[0]~0_combout ),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_31),
	.prn(vcc));
defparam \MonDReg[31] .is_wysiwyg = "true";
defparam \MonDReg[31] .power_up = "low";

dffeas \MonDReg[11] (
	.clk(clk_clk),
	.d(jdo_14),
	.asdata(q_a_11),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\MonDReg[0]~1_combout ),
	.sload(\MonDReg[0]~0_combout ),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_11),
	.prn(vcc));
defparam \MonDReg[11] .is_wysiwyg = "true";
defparam \MonDReg[11] .power_up = "low";

dffeas \MonDReg[10] (
	.clk(clk_clk),
	.d(jdo_13),
	.asdata(q_a_10),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\MonDReg[0]~1_combout ),
	.sload(\MonDReg[0]~0_combout ),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_10),
	.prn(vcc));
defparam \MonDReg[10] .is_wysiwyg = "true";
defparam \MonDReg[10] .power_up = "low";

dffeas \MonDReg[9] (
	.clk(clk_clk),
	.d(jdo_12),
	.asdata(q_a_9),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\MonDReg[0]~1_combout ),
	.sload(\MonDReg[0]~0_combout ),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_9),
	.prn(vcc));
defparam \MonDReg[9] .is_wysiwyg = "true";
defparam \MonDReg[9] .power_up = "low";

dffeas waitrequest(
	.clk(clk_clk),
	.d(\waitrequest~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(waitrequest1),
	.prn(vcc));
defparam waitrequest.is_wysiwyg = "true";
defparam waitrequest.power_up = "low";

dffeas \MonDReg[0] (
	.clk(clk_clk),
	.d(\MonDReg~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_0),
	.prn(vcc));
defparam \MonDReg[0] .is_wysiwyg = "true";
defparam \MonDReg[0] .power_up = "low";

dffeas \MonDReg[1] (
	.clk(clk_clk),
	.d(\MonDReg~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_1),
	.prn(vcc));
defparam \MonDReg[1] .is_wysiwyg = "true";
defparam \MonDReg[1] .power_up = "low";

dffeas \MonDReg[3] (
	.clk(clk_clk),
	.d(\MonDReg~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_3),
	.prn(vcc));
defparam \MonDReg[3] .is_wysiwyg = "true";
defparam \MonDReg[3] .power_up = "low";

dffeas \MonDReg[18] (
	.clk(clk_clk),
	.d(\MonDReg~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_18),
	.prn(vcc));
defparam \MonDReg[18] .is_wysiwyg = "true";
defparam \MonDReg[18] .power_up = "low";

dffeas \MonDReg[4] (
	.clk(clk_clk),
	.d(\MonDReg~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_4),
	.prn(vcc));
defparam \MonDReg[4] .is_wysiwyg = "true";
defparam \MonDReg[4] .power_up = "low";

dffeas \MonDReg[8] (
	.clk(clk_clk),
	.d(\MonDReg~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_8),
	.prn(vcc));
defparam \MonDReg[8] .is_wysiwyg = "true";
defparam \MonDReg[8] .power_up = "low";

dffeas \MonDReg[5] (
	.clk(clk_clk),
	.d(\MonDReg~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_5),
	.prn(vcc));
defparam \MonDReg[5] .is_wysiwyg = "true";
defparam \MonDReg[5] .power_up = "low";

dffeas \MonDReg[29] (
	.clk(clk_clk),
	.d(\MonDReg~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_29),
	.prn(vcc));
defparam \MonDReg[29] .is_wysiwyg = "true";
defparam \MonDReg[29] .power_up = "low";

dffeas \MonDReg[12] (
	.clk(clk_clk),
	.d(\MonDReg~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~2_combout ),
	.q(MonDReg_12),
	.prn(vcc));
defparam \MonDReg[12] .is_wysiwyg = "true";
defparam \MonDReg[12] .power_up = "low";

dffeas \MonDReg[15] (
	.clk(clk_clk),
	.d(\MonDReg~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!take_no_action_ocimem_a),
	.q(MonDReg_15),
	.prn(vcc));
defparam \MonDReg[15] .is_wysiwyg = "true";
defparam \MonDReg[15] .power_up = "low";

cyclonev_lcell_comb \Add0~1_wirecell (
	.dataa(!\Add0~1_sumout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~1_wirecell_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~1_wirecell .extended_lut = "off";
defparam \Add0~1_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \Add0~1_wirecell .shared_arith = "off";

dffeas \MonAReg[10] (
	.clk(clk_clk),
	.d(\Add0~1_wirecell_combout ),
	.asdata(jdo_17),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(take_action_ocimem_a1),
	.ena(take_action_ocimem_a),
	.q(\MonAReg[10]~q ),
	.prn(vcc));
defparam \MonAReg[10] .is_wysiwyg = "true";
defparam \MonAReg[10] .power_up = "low";

cyclonev_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\MonAReg[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout());
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h00000000000000FF;
defparam \Add0~9 .shared_arith = "off";

dffeas \MonAReg[2] (
	.clk(clk_clk),
	.d(\Add0~9_sumout ),
	.asdata(jdo_26),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(take_action_ocimem_a1),
	.ena(take_action_ocimem_a),
	.q(\MonAReg[2]~q ),
	.prn(vcc));
defparam \MonAReg[2] .is_wysiwyg = "true";
defparam \MonAReg[2] .power_up = "low";

cyclonev_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\MonAReg[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout());
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h00000000000000FF;
defparam \Add0~5 .shared_arith = "off";

dffeas \MonAReg[3] (
	.clk(clk_clk),
	.d(\Add0~5_sumout ),
	.asdata(jdo_27),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(take_action_ocimem_a1),
	.ena(take_action_ocimem_a),
	.q(\MonAReg[3]~q ),
	.prn(vcc));
defparam \MonAReg[3] .is_wysiwyg = "true";
defparam \MonAReg[3] .power_up = "low";

cyclonev_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\MonAReg[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout());
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h00000000000000FF;
defparam \Add0~13 .shared_arith = "off";

dffeas \MonAReg[4] (
	.clk(clk_clk),
	.d(\Add0~13_sumout ),
	.asdata(jdo_28),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(take_action_ocimem_a1),
	.ena(take_action_ocimem_a),
	.q(\MonAReg[4]~q ),
	.prn(vcc));
defparam \MonAReg[4] .is_wysiwyg = "true";
defparam \MonAReg[4] .power_up = "low";

cyclonev_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\MonAReg[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout());
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h00000000000000FF;
defparam \Add0~21 .shared_arith = "off";

dffeas \MonAReg[5] (
	.clk(clk_clk),
	.d(\Add0~21_sumout ),
	.asdata(jdo_29),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(take_action_ocimem_a1),
	.ena(take_action_ocimem_a),
	.q(\MonAReg[5]~q ),
	.prn(vcc));
defparam \MonAReg[5] .is_wysiwyg = "true";
defparam \MonAReg[5] .power_up = "low";

cyclonev_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\MonAReg[6]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout());
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h00000000000000FF;
defparam \Add0~25 .shared_arith = "off";

dffeas \MonAReg[6] (
	.clk(clk_clk),
	.d(\Add0~25_sumout ),
	.asdata(jdo_30),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(take_action_ocimem_a1),
	.ena(take_action_ocimem_a),
	.q(\MonAReg[6]~q ),
	.prn(vcc));
defparam \MonAReg[6] .is_wysiwyg = "true";
defparam \MonAReg[6] .power_up = "low";

cyclonev_lcell_comb \Add0~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\MonAReg[7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~29_sumout ),
	.cout(\Add0~30 ),
	.shareout());
defparam \Add0~29 .extended_lut = "off";
defparam \Add0~29 .lut_mask = 64'h00000000000000FF;
defparam \Add0~29 .shared_arith = "off";

dffeas \MonAReg[7] (
	.clk(clk_clk),
	.d(\Add0~29_sumout ),
	.asdata(jdo_31),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(take_action_ocimem_a1),
	.ena(take_action_ocimem_a),
	.q(\MonAReg[7]~q ),
	.prn(vcc));
defparam \MonAReg[7] .is_wysiwyg = "true";
defparam \MonAReg[7] .power_up = "low";

cyclonev_lcell_comb \Add0~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\MonAReg[8]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~33_sumout ),
	.cout(\Add0~34 ),
	.shareout());
defparam \Add0~33 .extended_lut = "off";
defparam \Add0~33 .lut_mask = 64'h00000000000000FF;
defparam \Add0~33 .shared_arith = "off";

dffeas \MonAReg[8] (
	.clk(clk_clk),
	.d(\Add0~33_sumout ),
	.asdata(jdo_32),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(take_action_ocimem_a1),
	.ena(take_action_ocimem_a),
	.q(\MonAReg[8]~q ),
	.prn(vcc));
defparam \MonAReg[8] .is_wysiwyg = "true";
defparam \MonAReg[8] .power_up = "low";

cyclonev_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\MonAReg[9]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout());
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h00000000000000FF;
defparam \Add0~17 .shared_arith = "off";

dffeas \MonAReg[9] (
	.clk(clk_clk),
	.d(\Add0~17_sumout ),
	.asdata(jdo_33),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(take_action_ocimem_a1),
	.ena(take_action_ocimem_a),
	.q(\MonAReg[9]~q ),
	.prn(vcc));
defparam \MonAReg[9] .is_wysiwyg = "true";
defparam \MonAReg[9] .power_up = "low";

cyclonev_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\MonAReg[10]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h00000000000000FF;
defparam \Add0~1 .shared_arith = "off";

cyclonev_lcell_comb \jtag_ram_rd~0 (
	.dataa(!jdo_34),
	.datab(!take_no_action_ocimem_a),
	.datac(!jdo_17),
	.datad(!\Add0~1_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\jtag_ram_rd~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \jtag_ram_rd~0 .extended_lut = "off";
defparam \jtag_ram_rd~0 .lut_mask = 64'hB1FFB1FFB1FFB1FF;
defparam \jtag_ram_rd~0 .shared_arith = "off";

cyclonev_lcell_comb \MonDReg[0]~0 (
	.dataa(!jdo_35),
	.datab(!take_action_ocimem_a),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\MonDReg[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \MonDReg[0]~0 .extended_lut = "off";
defparam \MonDReg[0]~0 .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \MonDReg[0]~0 .shared_arith = "off";

dffeas jtag_ram_rd(
	.clk(clk_clk),
	.d(\jtag_ram_rd~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~0_combout ),
	.q(\jtag_ram_rd~q ),
	.prn(vcc));
defparam jtag_ram_rd.is_wysiwyg = "true";
defparam jtag_ram_rd.power_up = "low";

dffeas jtag_ram_rd_d1(
	.clk(clk_clk),
	.d(\jtag_ram_rd~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\jtag_ram_rd_d1~q ),
	.prn(vcc));
defparam jtag_ram_rd_d1.is_wysiwyg = "true";
defparam jtag_ram_rd_d1.power_up = "low";

cyclonev_lcell_comb \MonDReg[0]~1 (
	.dataa(!\jtag_ram_rd_d1~q ),
	.datab(!\MonDReg[0]~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\MonDReg[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \MonDReg[0]~1 .extended_lut = "off";
defparam \MonDReg[0]~1 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \MonDReg[0]~1 .shared_arith = "off";

dffeas jtag_rd(
	.clk(clk_clk),
	.d(take_no_action_ocimem_a),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~0_combout ),
	.q(\jtag_rd~q ),
	.prn(vcc));
defparam jtag_rd.is_wysiwyg = "true";
defparam jtag_rd.power_up = "low";

dffeas jtag_rd_d1(
	.clk(clk_clk),
	.d(\jtag_rd~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\jtag_rd_d1~q ),
	.prn(vcc));
defparam jtag_rd_d1.is_wysiwyg = "true";
defparam jtag_rd_d1.power_up = "low";

cyclonev_lcell_comb \MonDReg[0]~2 (
	.dataa(!jdo_35),
	.datab(!take_action_ocimem_a),
	.datac(!\jtag_rd_d1~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\MonDReg[0]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \MonDReg[0]~2 .extended_lut = "off";
defparam \MonDReg[0]~2 .lut_mask = 64'h4747474747474747;
defparam \MonDReg[0]~2 .shared_arith = "off";

cyclonev_lcell_comb \jtag_ram_access~0 (
	.dataa(!jdo_34),
	.datab(!jdo_35),
	.datac(!take_action_ocimem_a),
	.datad(!jdo_17),
	.datae(!\Add0~1_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\jtag_ram_access~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \jtag_ram_access~0 .extended_lut = "off";
defparam \jtag_ram_access~0 .lut_mask = 64'hFF6FFFFFFF6FFFFF;
defparam \jtag_ram_access~0 .shared_arith = "off";

dffeas jtag_ram_access(
	.clk(clk_clk),
	.d(\jtag_ram_access~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\jtag_ram_access~q ),
	.prn(vcc));
defparam jtag_ram_access.is_wysiwyg = "true";
defparam jtag_ram_access.power_up = "low";

cyclonev_lcell_comb \waitrequest~0 (
	.dataa(!address_8),
	.datab(!\jtag_ram_access~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\waitrequest~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \waitrequest~0 .extended_lut = "off";
defparam \waitrequest~0 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \waitrequest~0 .shared_arith = "off";

cyclonev_lcell_comb \avalon_ociram_readdata_ready~0 (
	.dataa(!waitrequest1),
	.datab(!write),
	.datac(!\waitrequest~0_combout ),
	.datad(!read),
	.datae(!\avalon_ociram_readdata_ready~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\avalon_ociram_readdata_ready~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \avalon_ociram_readdata_ready~0 .extended_lut = "off";
defparam \avalon_ociram_readdata_ready~0 .lut_mask = 64'hD1FFFFFFD1FFFFFF;
defparam \avalon_ociram_readdata_ready~0 .shared_arith = "off";

dffeas avalon_ociram_readdata_ready(
	.clk(clk_clk),
	.d(\avalon_ociram_readdata_ready~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\avalon_ociram_readdata_ready~q ),
	.prn(vcc));
defparam avalon_ociram_readdata_ready.is_wysiwyg = "true";
defparam avalon_ociram_readdata_ready.power_up = "low";

cyclonev_lcell_comb \waitrequest~1 (
	.dataa(!waitrequest1),
	.datab(!write),
	.datac(!\waitrequest~0_combout ),
	.datad(!read),
	.datae(!\avalon_ociram_readdata_ready~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\waitrequest~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \waitrequest~1 .extended_lut = "off";
defparam \waitrequest~1 .lut_mask = 64'hFFFFBF8FFFFFBF8F;
defparam \waitrequest~1 .shared_arith = "off";

cyclonev_lcell_comb \MonDReg~15 (
	.dataa(!\MonAReg[4]~q ),
	.datab(!\MonAReg[2]~q ),
	.datac(!\jtag_ram_rd_d1~q ),
	.datad(!\MonAReg[3]~q ),
	.datae(!\MonDReg[0]~0_combout ),
	.dataf(!q_a_0),
	.datag(!jdo_3),
	.cin(gnd),
	.sharein(gnd),
	.combout(\MonDReg~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \MonDReg~15 .extended_lut = "on";
defparam \MonDReg~15 .lut_mask = 64'hF6FF96FFF6FF96FF;
defparam \MonDReg~15 .shared_arith = "off";

cyclonev_lcell_comb \Equal0~0 (
	.dataa(!\MonAReg[3]~q ),
	.datab(!\MonAReg[2]~q ),
	.datac(!\MonAReg[4]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~0 .extended_lut = "off";
defparam \Equal0~0 .lut_mask = 64'hEFEFEFEFEFEFEFEF;
defparam \Equal0~0 .shared_arith = "off";

cyclonev_lcell_comb \MonDReg~3 (
	.dataa(!\jtag_ram_rd_d1~q ),
	.datab(!\MonDReg[0]~0_combout ),
	.datac(!\Equal0~0_combout ),
	.datad(!jdo_4),
	.datae(!q_a_1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\MonDReg~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \MonDReg~3 .extended_lut = "off";
defparam \MonDReg~3 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \MonDReg~3 .shared_arith = "off";

cyclonev_lcell_comb \MonDReg~4 (
	.dataa(!\jtag_ram_rd_d1~q ),
	.datab(!\MonDReg[0]~0_combout ),
	.datac(!\Equal0~0_combout ),
	.datad(!q_a_3),
	.datae(!jdo_6),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\MonDReg~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \MonDReg~4 .extended_lut = "off";
defparam \MonDReg~4 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \MonDReg~4 .shared_arith = "off";

cyclonev_lcell_comb \MonDReg~12 (
	.dataa(!\MonAReg[2]~q ),
	.datab(!\MonAReg[4]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\MonDReg~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \MonDReg~12 .extended_lut = "off";
defparam \MonDReg~12 .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \MonDReg~12 .shared_arith = "off";

cyclonev_lcell_comb \MonDReg~5 (
	.dataa(!jdo_21),
	.datab(!\MonDReg[0]~0_combout ),
	.datac(!\MonAReg[3]~q ),
	.datad(!\jtag_ram_rd_d1~q ),
	.datae(!q_a_18),
	.dataf(!\MonDReg~12_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\MonDReg~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \MonDReg~5 .extended_lut = "off";
defparam \MonDReg~5 .lut_mask = 64'h7FDFFFFFFFFFFFFF;
defparam \MonDReg~5 .shared_arith = "off";

cyclonev_lcell_comb \MonDReg~6 (
	.dataa(!\MonAReg[3]~q ),
	.datab(!\MonAReg[2]~q ),
	.datac(!\MonAReg[4]~q ),
	.datad(!\jtag_ram_rd_d1~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\MonDReg~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \MonDReg~6 .extended_lut = "off";
defparam \MonDReg~6 .lut_mask = 64'hFFFBFFFBFFFBFFFB;
defparam \MonDReg~6 .shared_arith = "off";

cyclonev_lcell_comb \MonDReg~7 (
	.dataa(!\jtag_ram_rd_d1~q ),
	.datab(!\MonDReg[0]~0_combout ),
	.datac(!q_a_4),
	.datad(!jdo_7),
	.datae(!\MonDReg~6_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\MonDReg~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \MonDReg~7 .extended_lut = "off";
defparam \MonDReg~7 .lut_mask = 64'h47FFFFFF47FFFFFF;
defparam \MonDReg~7 .shared_arith = "off";

cyclonev_lcell_comb \MonDReg~14 (
	.dataa(!\MonDReg[0]~0_combout ),
	.datab(!\jtag_ram_rd_d1~q ),
	.datac(!\MonAReg[4]~q ),
	.datad(!\MonAReg[2]~q ),
	.datae(!q_a_8),
	.dataf(!jdo_11),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\MonDReg~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \MonDReg~14 .extended_lut = "off";
defparam \MonDReg~14 .lut_mask = 64'hF6FFFFFFFFFFFFFF;
defparam \MonDReg~14 .shared_arith = "off";

cyclonev_lcell_comb \Equal0~1 (
	.dataa(!\MonAReg[3]~q ),
	.datab(!\MonAReg[2]~q ),
	.datac(!\MonAReg[4]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~1 .extended_lut = "off";
defparam \Equal0~1 .lut_mask = 64'hFEFEFEFEFEFEFEFE;
defparam \Equal0~1 .shared_arith = "off";

cyclonev_lcell_comb \MonDReg~8 (
	.dataa(!\Equal0~1_combout ),
	.datab(!\jtag_ram_rd_d1~q ),
	.datac(!\MonDReg[0]~0_combout ),
	.datad(!q_a_5),
	.datae(!jdo_8),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\MonDReg~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \MonDReg~8 .extended_lut = "off";
defparam \MonDReg~8 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \MonDReg~8 .shared_arith = "off";

cyclonev_lcell_comb \MonDReg~9 (
	.dataa(!\jtag_ram_rd_d1~q ),
	.datab(!\MonDReg[0]~0_combout ),
	.datac(!\Equal0~0_combout ),
	.datad(!jdo_32),
	.datae(!q_a_29),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\MonDReg~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \MonDReg~9 .extended_lut = "off";
defparam \MonDReg~9 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \MonDReg~9 .shared_arith = "off";

cyclonev_lcell_comb \MonDReg~10 (
	.dataa(!\jtag_ram_rd_d1~q ),
	.datab(!\MonDReg[0]~0_combout ),
	.datac(!q_a_12),
	.datad(!\MonDReg~6_combout ),
	.datae(!jdo_15),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\MonDReg~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \MonDReg~10 .extended_lut = "off";
defparam \MonDReg~10 .lut_mask = 64'h47FFFFFF47FFFFFF;
defparam \MonDReg~10 .shared_arith = "off";

cyclonev_lcell_comb \MonDReg~13 (
	.dataa(!\jtag_rd_d1~q ),
	.datab(!MonDReg_15),
	.datac(!\MonAReg[3]~q ),
	.datad(!\MonAReg[2]~q ),
	.datae(!\MonAReg[4]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\MonDReg~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \MonDReg~13 .extended_lut = "off";
defparam \MonDReg~13 .lut_mask = 64'hFBF7F7FBFBF7F7FB;
defparam \MonDReg~13 .shared_arith = "off";

cyclonev_lcell_comb \MonDReg~11 (
	.dataa(!\MonDReg[0]~0_combout ),
	.datab(!\jtag_rd_d1~q ),
	.datac(!jdo_18),
	.datad(!\jtag_ram_rd_d1~q ),
	.datae(!q_a_15),
	.dataf(!\MonDReg~13_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\MonDReg~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \MonDReg~11 .extended_lut = "off";
defparam \MonDReg~11 .lut_mask = 64'h9F6FFFFFFFFFFFFF;
defparam \MonDReg~11 .shared_arith = "off";

endmodule

module processor_processor_cpu_ociram_sp_ram_module (
	q_a_0,
	q_a_1,
	q_a_2,
	q_a_16,
	q_a_8,
	q_a_24,
	q_a_20,
	q_a_19,
	q_a_5,
	q_a_21,
	q_a_13,
	q_a_29,
	q_a_4,
	q_a_12,
	q_a_28,
	q_a_6,
	q_a_22,
	q_a_14,
	q_a_30,
	q_a_7,
	q_a_23,
	q_a_15,
	q_a_31,
	q_a_11,
	q_a_27,
	q_a_10,
	q_a_26,
	q_a_25,
	q_a_9,
	q_a_3,
	q_a_18,
	q_a_17,
	ociram_wr_en,
	ociram_reset_req,
	ociram_wr_data_0,
	ociram_addr_0,
	ociram_addr_1,
	ociram_addr_2,
	ociram_addr_3,
	ociram_addr_4,
	ociram_addr_5,
	ociram_addr_6,
	ociram_addr_7,
	ociram_byteenable_0,
	ociram_wr_data_1,
	ociram_wr_data_2,
	ociram_wr_data_16,
	ociram_byteenable_2,
	ociram_wr_data_8,
	ociram_byteenable_1,
	ociram_wr_data_24,
	ociram_byteenable_3,
	ociram_wr_data_20,
	ociram_wr_data_19,
	ociram_wr_data_5,
	ociram_wr_data_21,
	ociram_wr_data_13,
	ociram_wr_data_29,
	ociram_wr_data_4,
	ociram_wr_data_12,
	ociram_wr_data_28,
	ociram_wr_data_6,
	ociram_wr_data_22,
	ociram_wr_data_14,
	ociram_wr_data_30,
	ociram_wr_data_7,
	ociram_wr_data_23,
	ociram_wr_data_15,
	ociram_wr_data_31,
	ociram_wr_data_11,
	ociram_wr_data_27,
	ociram_wr_data_10,
	ociram_wr_data_26,
	ociram_wr_data_25,
	ociram_wr_data_9,
	ociram_wr_data_3,
	ociram_wr_data_18,
	ociram_wr_data_17,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	q_a_0;
output 	q_a_1;
output 	q_a_2;
output 	q_a_16;
output 	q_a_8;
output 	q_a_24;
output 	q_a_20;
output 	q_a_19;
output 	q_a_5;
output 	q_a_21;
output 	q_a_13;
output 	q_a_29;
output 	q_a_4;
output 	q_a_12;
output 	q_a_28;
output 	q_a_6;
output 	q_a_22;
output 	q_a_14;
output 	q_a_30;
output 	q_a_7;
output 	q_a_23;
output 	q_a_15;
output 	q_a_31;
output 	q_a_11;
output 	q_a_27;
output 	q_a_10;
output 	q_a_26;
output 	q_a_25;
output 	q_a_9;
output 	q_a_3;
output 	q_a_18;
output 	q_a_17;
input 	ociram_wr_en;
input 	ociram_reset_req;
input 	ociram_wr_data_0;
input 	ociram_addr_0;
input 	ociram_addr_1;
input 	ociram_addr_2;
input 	ociram_addr_3;
input 	ociram_addr_4;
input 	ociram_addr_5;
input 	ociram_addr_6;
input 	ociram_addr_7;
input 	ociram_byteenable_0;
input 	ociram_wr_data_1;
input 	ociram_wr_data_2;
input 	ociram_wr_data_16;
input 	ociram_byteenable_2;
input 	ociram_wr_data_8;
input 	ociram_byteenable_1;
input 	ociram_wr_data_24;
input 	ociram_byteenable_3;
input 	ociram_wr_data_20;
input 	ociram_wr_data_19;
input 	ociram_wr_data_5;
input 	ociram_wr_data_21;
input 	ociram_wr_data_13;
input 	ociram_wr_data_29;
input 	ociram_wr_data_4;
input 	ociram_wr_data_12;
input 	ociram_wr_data_28;
input 	ociram_wr_data_6;
input 	ociram_wr_data_22;
input 	ociram_wr_data_14;
input 	ociram_wr_data_30;
input 	ociram_wr_data_7;
input 	ociram_wr_data_23;
input 	ociram_wr_data_15;
input 	ociram_wr_data_31;
input 	ociram_wr_data_11;
input 	ociram_wr_data_27;
input 	ociram_wr_data_10;
input 	ociram_wr_data_26;
input 	ociram_wr_data_25;
input 	ociram_wr_data_9;
input 	ociram_wr_data_3;
input 	ociram_wr_data_18;
input 	ociram_wr_data_17;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



processor_altsyncram_3 the_altsyncram(
	.q_a({q_a_31,q_a_30,q_a_29,q_a_28,q_a_27,q_a_26,q_a_25,q_a_24,q_a_23,q_a_22,q_a_21,q_a_20,q_a_19,q_a_18,q_a_17,q_a_16,q_a_15,q_a_14,q_a_13,q_a_12,q_a_11,q_a_10,q_a_9,q_a_8,q_a_7,q_a_6,q_a_5,q_a_4,q_a_3,q_a_2,q_a_1,q_a_0}),
	.wren_a(ociram_wr_en),
	.clocken0(ociram_reset_req),
	.data_a({ociram_wr_data_31,ociram_wr_data_30,ociram_wr_data_29,ociram_wr_data_28,ociram_wr_data_27,ociram_wr_data_26,ociram_wr_data_25,ociram_wr_data_24,ociram_wr_data_23,ociram_wr_data_22,ociram_wr_data_21,ociram_wr_data_20,ociram_wr_data_19,ociram_wr_data_18,ociram_wr_data_17,
ociram_wr_data_16,ociram_wr_data_15,ociram_wr_data_14,ociram_wr_data_13,ociram_wr_data_12,ociram_wr_data_11,ociram_wr_data_10,ociram_wr_data_9,ociram_wr_data_8,ociram_wr_data_7,ociram_wr_data_6,ociram_wr_data_5,ociram_wr_data_4,ociram_wr_data_3,ociram_wr_data_2,
ociram_wr_data_1,ociram_wr_data_0}),
	.address_a({gnd,gnd,gnd,gnd,gnd,ociram_addr_7,ociram_addr_6,ociram_addr_5,ociram_addr_4,ociram_addr_3,ociram_addr_2,ociram_addr_1,ociram_addr_0}),
	.byteena_a({ociram_byteenable_3,ociram_byteenable_2,ociram_byteenable_1,ociram_byteenable_0}),
	.clock0(clk_clk));

endmodule

module processor_altsyncram_3 (
	q_a,
	wren_a,
	clocken0,
	data_a,
	address_a,
	byteena_a,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[31:0] q_a;
input 	wren_a;
input 	clocken0;
input 	[31:0] data_a;
input 	[12:0] address_a;
input 	[3:0] byteena_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



processor_altsyncram_4qe1 auto_generated(
	.q_a({q_a[31],q_a[30],q_a[29],q_a[28],q_a[27],q_a[26],q_a[25],q_a[24],q_a[23],q_a[22],q_a[21],q_a[20],q_a[19],q_a[18],q_a[17],q_a[16],q_a[15],q_a[14],q_a[13],q_a[12],q_a[11],q_a[10],q_a[9],q_a[8],q_a[7],q_a[6],q_a[5],q_a[4],q_a[3],q_a[2],q_a[1],q_a[0]}),
	.wren_a(wren_a),
	.clocken0(clocken0),
	.data_a({data_a[31],data_a[30],data_a[29],data_a[28],data_a[27],data_a[26],data_a[25],data_a[24],data_a[23],data_a[22],data_a[21],data_a[20],data_a[19],data_a[18],data_a[17],data_a[16],data_a[15],data_a[14],data_a[13],data_a[12],data_a[11],data_a[10],data_a[9],data_a[8],data_a[7],data_a[6],data_a[5],data_a[4],data_a[3],data_a[2],data_a[1],data_a[0]}),
	.address_a({address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.byteena_a({byteena_a[3],byteena_a[2],byteena_a[1],byteena_a[0]}),
	.clock0(clock0));

endmodule

module processor_altsyncram_4qe1 (
	q_a,
	wren_a,
	clocken0,
	data_a,
	address_a,
	byteena_a,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[31:0] q_a;
input 	wren_a;
input 	clocken0;
input 	[31:0] data_a;
input 	[7:0] address_a;
input 	[3:0] byteena_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a0_PORTADATAOUT_bus;
wire [143:0] ram_block1a1_PORTADATAOUT_bus;
wire [143:0] ram_block1a2_PORTADATAOUT_bus;
wire [143:0] ram_block1a16_PORTADATAOUT_bus;
wire [143:0] ram_block1a8_PORTADATAOUT_bus;
wire [143:0] ram_block1a24_PORTADATAOUT_bus;
wire [143:0] ram_block1a20_PORTADATAOUT_bus;
wire [143:0] ram_block1a19_PORTADATAOUT_bus;
wire [143:0] ram_block1a5_PORTADATAOUT_bus;
wire [143:0] ram_block1a21_PORTADATAOUT_bus;
wire [143:0] ram_block1a13_PORTADATAOUT_bus;
wire [143:0] ram_block1a29_PORTADATAOUT_bus;
wire [143:0] ram_block1a4_PORTADATAOUT_bus;
wire [143:0] ram_block1a12_PORTADATAOUT_bus;
wire [143:0] ram_block1a28_PORTADATAOUT_bus;
wire [143:0] ram_block1a6_PORTADATAOUT_bus;
wire [143:0] ram_block1a22_PORTADATAOUT_bus;
wire [143:0] ram_block1a14_PORTADATAOUT_bus;
wire [143:0] ram_block1a30_PORTADATAOUT_bus;
wire [143:0] ram_block1a7_PORTADATAOUT_bus;
wire [143:0] ram_block1a23_PORTADATAOUT_bus;
wire [143:0] ram_block1a15_PORTADATAOUT_bus;
wire [143:0] ram_block1a31_PORTADATAOUT_bus;
wire [143:0] ram_block1a11_PORTADATAOUT_bus;
wire [143:0] ram_block1a27_PORTADATAOUT_bus;
wire [143:0] ram_block1a10_PORTADATAOUT_bus;
wire [143:0] ram_block1a26_PORTADATAOUT_bus;
wire [143:0] ram_block1a25_PORTADATAOUT_bus;
wire [143:0] ram_block1a9_PORTADATAOUT_bus;
wire [143:0] ram_block1a3_PORTADATAOUT_bus;
wire [143:0] ram_block1a18_PORTADATAOUT_bus;
wire [143:0] ram_block1a17_PORTADATAOUT_bus;

assign q_a[0] = ram_block1a0_PORTADATAOUT_bus[0];

assign q_a[1] = ram_block1a1_PORTADATAOUT_bus[0];

assign q_a[2] = ram_block1a2_PORTADATAOUT_bus[0];

assign q_a[16] = ram_block1a16_PORTADATAOUT_bus[0];

assign q_a[8] = ram_block1a8_PORTADATAOUT_bus[0];

assign q_a[24] = ram_block1a24_PORTADATAOUT_bus[0];

assign q_a[20] = ram_block1a20_PORTADATAOUT_bus[0];

assign q_a[19] = ram_block1a19_PORTADATAOUT_bus[0];

assign q_a[5] = ram_block1a5_PORTADATAOUT_bus[0];

assign q_a[21] = ram_block1a21_PORTADATAOUT_bus[0];

assign q_a[13] = ram_block1a13_PORTADATAOUT_bus[0];

assign q_a[29] = ram_block1a29_PORTADATAOUT_bus[0];

assign q_a[4] = ram_block1a4_PORTADATAOUT_bus[0];

assign q_a[12] = ram_block1a12_PORTADATAOUT_bus[0];

assign q_a[28] = ram_block1a28_PORTADATAOUT_bus[0];

assign q_a[6] = ram_block1a6_PORTADATAOUT_bus[0];

assign q_a[22] = ram_block1a22_PORTADATAOUT_bus[0];

assign q_a[14] = ram_block1a14_PORTADATAOUT_bus[0];

assign q_a[30] = ram_block1a30_PORTADATAOUT_bus[0];

assign q_a[7] = ram_block1a7_PORTADATAOUT_bus[0];

assign q_a[23] = ram_block1a23_PORTADATAOUT_bus[0];

assign q_a[15] = ram_block1a15_PORTADATAOUT_bus[0];

assign q_a[31] = ram_block1a31_PORTADATAOUT_bus[0];

assign q_a[11] = ram_block1a11_PORTADATAOUT_bus[0];

assign q_a[27] = ram_block1a27_PORTADATAOUT_bus[0];

assign q_a[10] = ram_block1a10_PORTADATAOUT_bus[0];

assign q_a[26] = ram_block1a26_PORTADATAOUT_bus[0];

assign q_a[25] = ram_block1a25_PORTADATAOUT_bus[0];

assign q_a[9] = ram_block1a9_PORTADATAOUT_bus[0];

assign q_a[3] = ram_block1a3_PORTADATAOUT_bus[0];

assign q_a[18] = ram_block1a18_PORTADATAOUT_bus[0];

assign q_a[17] = ram_block1a17_PORTADATAOUT_bus[0];

cyclonev_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a0_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.clk0_input_clock_enable = "ena0";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.init_file = "processor_cpu_ociram_default_contents.mif";
defparam ram_block1a0.init_file_layout = "port_a";
defparam ram_block1a0.logical_ram_name = "processor_cpu:cpu|processor_cpu_nios2_oci:the_processor_cpu_nios2_oci|processor_cpu_nios2_ocimem:the_processor_cpu_nios2_ocimem|processor_cpu_ociram_sp_ram_module:processor_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_4qe1:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.operation_mode = "single_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 8;
defparam ram_block1a0.port_a_byte_enable_mask_width = 1;
defparam ram_block1a0.port_a_byte_size = 1;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 255;
defparam ram_block1a0.port_a_logical_ram_depth = 256;
defparam ram_block1a0.port_a_logical_ram_width = 32;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.ram_block_type = "auto";
defparam ram_block1a0.mem_init0 = "F082E980277062912CB244CFD084FC8EC49C6B4F28A560069238B1A3C7D5FBB6";

cyclonev_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a1_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a1.clk0_core_clock_enable = "ena0";
defparam ram_block1a1.clk0_input_clock_enable = "ena0";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.init_file = "processor_cpu_ociram_default_contents.mif";
defparam ram_block1a1.init_file_layout = "port_a";
defparam ram_block1a1.logical_ram_name = "processor_cpu:cpu|processor_cpu_nios2_oci:the_processor_cpu_nios2_oci|processor_cpu_nios2_ocimem:the_processor_cpu_nios2_ocimem|processor_cpu_ociram_sp_ram_module:processor_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_4qe1:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.operation_mode = "single_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 8;
defparam ram_block1a1.port_a_byte_enable_mask_width = 1;
defparam ram_block1a1.port_a_byte_size = 1;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 255;
defparam ram_block1a1.port_a_logical_ram_depth = 256;
defparam ram_block1a1.port_a_logical_ram_width = 32;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.ram_block_type = "auto";
defparam ram_block1a1.mem_init0 = "D79799D62A2EBCDE87554821870A4291446385CAE645D15F127F51099EE7FA77";

cyclonev_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a2_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a2.clk0_core_clock_enable = "ena0";
defparam ram_block1a2.clk0_input_clock_enable = "ena0";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.init_file = "processor_cpu_ociram_default_contents.mif";
defparam ram_block1a2.init_file_layout = "port_a";
defparam ram_block1a2.logical_ram_name = "processor_cpu:cpu|processor_cpu_nios2_oci:the_processor_cpu_nios2_oci|processor_cpu_nios2_ocimem:the_processor_cpu_nios2_ocimem|processor_cpu_ociram_sp_ram_module:processor_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_4qe1:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.operation_mode = "single_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 8;
defparam ram_block1a2.port_a_byte_enable_mask_width = 1;
defparam ram_block1a2.port_a_byte_size = 1;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 255;
defparam ram_block1a2.port_a_logical_ram_depth = 256;
defparam ram_block1a2.port_a_logical_ram_width = 32;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.ram_block_type = "auto";
defparam ram_block1a2.mem_init0 = "706E6722D5D1FDC707F573CF0D406D54B651FC97C911E5D3A44C8EF6E86E2CAE";

cyclonev_ram_block ram_block1a16(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a16_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a16.clk0_core_clock_enable = "ena0";
defparam ram_block1a16.clk0_input_clock_enable = "ena0";
defparam ram_block1a16.data_interleave_offset_in_bits = 1;
defparam ram_block1a16.data_interleave_width_in_bits = 1;
defparam ram_block1a16.init_file = "processor_cpu_ociram_default_contents.mif";
defparam ram_block1a16.init_file_layout = "port_a";
defparam ram_block1a16.logical_ram_name = "processor_cpu:cpu|processor_cpu_nios2_oci:the_processor_cpu_nios2_oci|processor_cpu_nios2_ocimem:the_processor_cpu_nios2_ocimem|processor_cpu_ociram_sp_ram_module:processor_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_4qe1:auto_generated|ALTSYNCRAM";
defparam ram_block1a16.operation_mode = "single_port";
defparam ram_block1a16.port_a_address_clear = "none";
defparam ram_block1a16.port_a_address_width = 8;
defparam ram_block1a16.port_a_byte_enable_mask_width = 1;
defparam ram_block1a16.port_a_byte_size = 1;
defparam ram_block1a16.port_a_data_out_clear = "none";
defparam ram_block1a16.port_a_data_out_clock = "none";
defparam ram_block1a16.port_a_data_width = 1;
defparam ram_block1a16.port_a_first_address = 0;
defparam ram_block1a16.port_a_first_bit_number = 16;
defparam ram_block1a16.port_a_last_address = 255;
defparam ram_block1a16.port_a_logical_ram_depth = 256;
defparam ram_block1a16.port_a_logical_ram_width = 32;
defparam ram_block1a16.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a16.ram_block_type = "auto";
defparam ram_block1a16.mem_init0 = "A5D90182D0FEE54279153DC162279DA35E59C350C65ACE273B5053B17E638A67";

cyclonev_ram_block ram_block1a8(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a8_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a8.clk0_core_clock_enable = "ena0";
defparam ram_block1a8.clk0_input_clock_enable = "ena0";
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.init_file = "processor_cpu_ociram_default_contents.mif";
defparam ram_block1a8.init_file_layout = "port_a";
defparam ram_block1a8.logical_ram_name = "processor_cpu:cpu|processor_cpu_nios2_oci:the_processor_cpu_nios2_oci|processor_cpu_nios2_ocimem:the_processor_cpu_nios2_ocimem|processor_cpu_ociram_sp_ram_module:processor_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_4qe1:auto_generated|ALTSYNCRAM";
defparam ram_block1a8.operation_mode = "single_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 8;
defparam ram_block1a8.port_a_byte_enable_mask_width = 1;
defparam ram_block1a8.port_a_byte_size = 1;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 255;
defparam ram_block1a8.port_a_logical_ram_depth = 256;
defparam ram_block1a8.port_a_logical_ram_width = 32;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a8.ram_block_type = "auto";
defparam ram_block1a8.mem_init0 = "B4D77C1E3C88B38DC941C69776E33B1C652A6C84E88338640BBFAD3B06EF524E";

cyclonev_ram_block ram_block1a24(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[24]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a24_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a24.clk0_core_clock_enable = "ena0";
defparam ram_block1a24.clk0_input_clock_enable = "ena0";
defparam ram_block1a24.data_interleave_offset_in_bits = 1;
defparam ram_block1a24.data_interleave_width_in_bits = 1;
defparam ram_block1a24.init_file = "processor_cpu_ociram_default_contents.mif";
defparam ram_block1a24.init_file_layout = "port_a";
defparam ram_block1a24.logical_ram_name = "processor_cpu:cpu|processor_cpu_nios2_oci:the_processor_cpu_nios2_oci|processor_cpu_nios2_ocimem:the_processor_cpu_nios2_ocimem|processor_cpu_ociram_sp_ram_module:processor_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_4qe1:auto_generated|ALTSYNCRAM";
defparam ram_block1a24.operation_mode = "single_port";
defparam ram_block1a24.port_a_address_clear = "none";
defparam ram_block1a24.port_a_address_width = 8;
defparam ram_block1a24.port_a_byte_enable_mask_width = 1;
defparam ram_block1a24.port_a_byte_size = 1;
defparam ram_block1a24.port_a_data_out_clear = "none";
defparam ram_block1a24.port_a_data_out_clock = "none";
defparam ram_block1a24.port_a_data_width = 1;
defparam ram_block1a24.port_a_first_address = 0;
defparam ram_block1a24.port_a_first_bit_number = 24;
defparam ram_block1a24.port_a_last_address = 255;
defparam ram_block1a24.port_a_logical_ram_depth = 256;
defparam ram_block1a24.port_a_logical_ram_width = 32;
defparam ram_block1a24.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a24.ram_block_type = "auto";
defparam ram_block1a24.mem_init0 = "471DD74C4854A7C640358F5D02EF6605C204E43D414864177C2880AD9B4E5B41";

cyclonev_ram_block ram_block1a20(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[20]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a20_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a20.clk0_core_clock_enable = "ena0";
defparam ram_block1a20.clk0_input_clock_enable = "ena0";
defparam ram_block1a20.data_interleave_offset_in_bits = 1;
defparam ram_block1a20.data_interleave_width_in_bits = 1;
defparam ram_block1a20.init_file = "processor_cpu_ociram_default_contents.mif";
defparam ram_block1a20.init_file_layout = "port_a";
defparam ram_block1a20.logical_ram_name = "processor_cpu:cpu|processor_cpu_nios2_oci:the_processor_cpu_nios2_oci|processor_cpu_nios2_ocimem:the_processor_cpu_nios2_ocimem|processor_cpu_ociram_sp_ram_module:processor_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_4qe1:auto_generated|ALTSYNCRAM";
defparam ram_block1a20.operation_mode = "single_port";
defparam ram_block1a20.port_a_address_clear = "none";
defparam ram_block1a20.port_a_address_width = 8;
defparam ram_block1a20.port_a_byte_enable_mask_width = 1;
defparam ram_block1a20.port_a_byte_size = 1;
defparam ram_block1a20.port_a_data_out_clear = "none";
defparam ram_block1a20.port_a_data_out_clock = "none";
defparam ram_block1a20.port_a_data_width = 1;
defparam ram_block1a20.port_a_first_address = 0;
defparam ram_block1a20.port_a_first_bit_number = 20;
defparam ram_block1a20.port_a_last_address = 255;
defparam ram_block1a20.port_a_logical_ram_depth = 256;
defparam ram_block1a20.port_a_logical_ram_width = 32;
defparam ram_block1a20.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a20.ram_block_type = "auto";
defparam ram_block1a20.mem_init0 = "5CF4DC015DC4B93CAC73E3F541C878BD0279B1FC525FA32A7BD99A286AF85CDD";

cyclonev_ram_block ram_block1a19(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[19]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a19_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a19.clk0_core_clock_enable = "ena0";
defparam ram_block1a19.clk0_input_clock_enable = "ena0";
defparam ram_block1a19.data_interleave_offset_in_bits = 1;
defparam ram_block1a19.data_interleave_width_in_bits = 1;
defparam ram_block1a19.init_file = "processor_cpu_ociram_default_contents.mif";
defparam ram_block1a19.init_file_layout = "port_a";
defparam ram_block1a19.logical_ram_name = "processor_cpu:cpu|processor_cpu_nios2_oci:the_processor_cpu_nios2_oci|processor_cpu_nios2_ocimem:the_processor_cpu_nios2_ocimem|processor_cpu_ociram_sp_ram_module:processor_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_4qe1:auto_generated|ALTSYNCRAM";
defparam ram_block1a19.operation_mode = "single_port";
defparam ram_block1a19.port_a_address_clear = "none";
defparam ram_block1a19.port_a_address_width = 8;
defparam ram_block1a19.port_a_byte_enable_mask_width = 1;
defparam ram_block1a19.port_a_byte_size = 1;
defparam ram_block1a19.port_a_data_out_clear = "none";
defparam ram_block1a19.port_a_data_out_clock = "none";
defparam ram_block1a19.port_a_data_width = 1;
defparam ram_block1a19.port_a_first_address = 0;
defparam ram_block1a19.port_a_first_bit_number = 19;
defparam ram_block1a19.port_a_last_address = 255;
defparam ram_block1a19.port_a_logical_ram_depth = 256;
defparam ram_block1a19.port_a_logical_ram_width = 32;
defparam ram_block1a19.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a19.ram_block_type = "auto";
defparam ram_block1a19.mem_init0 = "360DDF4DBED01AA957F9DF48CA69E672F9EEDAFEAC738A5C72EF5CB7DDA7D30D";

cyclonev_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a5_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a5.clk0_core_clock_enable = "ena0";
defparam ram_block1a5.clk0_input_clock_enable = "ena0";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.init_file = "processor_cpu_ociram_default_contents.mif";
defparam ram_block1a5.init_file_layout = "port_a";
defparam ram_block1a5.logical_ram_name = "processor_cpu:cpu|processor_cpu_nios2_oci:the_processor_cpu_nios2_oci|processor_cpu_nios2_ocimem:the_processor_cpu_nios2_ocimem|processor_cpu_ociram_sp_ram_module:processor_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_4qe1:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.operation_mode = "single_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 8;
defparam ram_block1a5.port_a_byte_enable_mask_width = 1;
defparam ram_block1a5.port_a_byte_size = 1;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 255;
defparam ram_block1a5.port_a_logical_ram_depth = 256;
defparam ram_block1a5.port_a_logical_ram_width = 32;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.ram_block_type = "auto";
defparam ram_block1a5.mem_init0 = "56385C7763CD70C3C6A16547526E3BE75D897A6DE98AB7B6A2B89B3CBC1026F9";

cyclonev_ram_block ram_block1a21(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[21]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a21_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a21.clk0_core_clock_enable = "ena0";
defparam ram_block1a21.clk0_input_clock_enable = "ena0";
defparam ram_block1a21.data_interleave_offset_in_bits = 1;
defparam ram_block1a21.data_interleave_width_in_bits = 1;
defparam ram_block1a21.init_file = "processor_cpu_ociram_default_contents.mif";
defparam ram_block1a21.init_file_layout = "port_a";
defparam ram_block1a21.logical_ram_name = "processor_cpu:cpu|processor_cpu_nios2_oci:the_processor_cpu_nios2_oci|processor_cpu_nios2_ocimem:the_processor_cpu_nios2_ocimem|processor_cpu_ociram_sp_ram_module:processor_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_4qe1:auto_generated|ALTSYNCRAM";
defparam ram_block1a21.operation_mode = "single_port";
defparam ram_block1a21.port_a_address_clear = "none";
defparam ram_block1a21.port_a_address_width = 8;
defparam ram_block1a21.port_a_byte_enable_mask_width = 1;
defparam ram_block1a21.port_a_byte_size = 1;
defparam ram_block1a21.port_a_data_out_clear = "none";
defparam ram_block1a21.port_a_data_out_clock = "none";
defparam ram_block1a21.port_a_data_width = 1;
defparam ram_block1a21.port_a_first_address = 0;
defparam ram_block1a21.port_a_first_bit_number = 21;
defparam ram_block1a21.port_a_last_address = 255;
defparam ram_block1a21.port_a_logical_ram_depth = 256;
defparam ram_block1a21.port_a_logical_ram_width = 32;
defparam ram_block1a21.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a21.ram_block_type = "auto";
defparam ram_block1a21.mem_init0 = "B50B0604E542D1D67047F6548C867D78F987A48D04D1CA5CF25047175F2674EC";

cyclonev_ram_block ram_block1a13(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a13_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a13.clk0_core_clock_enable = "ena0";
defparam ram_block1a13.clk0_input_clock_enable = "ena0";
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.init_file = "processor_cpu_ociram_default_contents.mif";
defparam ram_block1a13.init_file_layout = "port_a";
defparam ram_block1a13.logical_ram_name = "processor_cpu:cpu|processor_cpu_nios2_oci:the_processor_cpu_nios2_oci|processor_cpu_nios2_ocimem:the_processor_cpu_nios2_ocimem|processor_cpu_ociram_sp_ram_module:processor_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_4qe1:auto_generated|ALTSYNCRAM";
defparam ram_block1a13.operation_mode = "single_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 8;
defparam ram_block1a13.port_a_byte_enable_mask_width = 1;
defparam ram_block1a13.port_a_byte_size = 1;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 255;
defparam ram_block1a13.port_a_logical_ram_depth = 256;
defparam ram_block1a13.port_a_logical_ram_width = 32;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a13.ram_block_type = "auto";
defparam ram_block1a13.mem_init0 = "D891C645AC0EC442B741340091FA518E10D334A5CC003D79760E04EBBDE9A522";

cyclonev_ram_block ram_block1a29(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[29]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a29_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a29.clk0_core_clock_enable = "ena0";
defparam ram_block1a29.clk0_input_clock_enable = "ena0";
defparam ram_block1a29.data_interleave_offset_in_bits = 1;
defparam ram_block1a29.data_interleave_width_in_bits = 1;
defparam ram_block1a29.init_file = "processor_cpu_ociram_default_contents.mif";
defparam ram_block1a29.init_file_layout = "port_a";
defparam ram_block1a29.logical_ram_name = "processor_cpu:cpu|processor_cpu_nios2_oci:the_processor_cpu_nios2_oci|processor_cpu_nios2_ocimem:the_processor_cpu_nios2_ocimem|processor_cpu_ociram_sp_ram_module:processor_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_4qe1:auto_generated|ALTSYNCRAM";
defparam ram_block1a29.operation_mode = "single_port";
defparam ram_block1a29.port_a_address_clear = "none";
defparam ram_block1a29.port_a_address_width = 8;
defparam ram_block1a29.port_a_byte_enable_mask_width = 1;
defparam ram_block1a29.port_a_byte_size = 1;
defparam ram_block1a29.port_a_data_out_clear = "none";
defparam ram_block1a29.port_a_data_out_clock = "none";
defparam ram_block1a29.port_a_data_width = 1;
defparam ram_block1a29.port_a_first_address = 0;
defparam ram_block1a29.port_a_first_bit_number = 29;
defparam ram_block1a29.port_a_last_address = 255;
defparam ram_block1a29.port_a_logical_ram_depth = 256;
defparam ram_block1a29.port_a_logical_ram_width = 32;
defparam ram_block1a29.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a29.ram_block_type = "auto";
defparam ram_block1a29.mem_init0 = "480F616A1CF268494538501BEFD54167C5679AB6979341F9D788674983C166D0";

cyclonev_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a4_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a4.clk0_core_clock_enable = "ena0";
defparam ram_block1a4.clk0_input_clock_enable = "ena0";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.init_file = "processor_cpu_ociram_default_contents.mif";
defparam ram_block1a4.init_file_layout = "port_a";
defparam ram_block1a4.logical_ram_name = "processor_cpu:cpu|processor_cpu_nios2_oci:the_processor_cpu_nios2_oci|processor_cpu_nios2_ocimem:the_processor_cpu_nios2_ocimem|processor_cpu_ociram_sp_ram_module:processor_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_4qe1:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.operation_mode = "single_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 8;
defparam ram_block1a4.port_a_byte_enable_mask_width = 1;
defparam ram_block1a4.port_a_byte_size = 1;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 255;
defparam ram_block1a4.port_a_logical_ram_depth = 256;
defparam ram_block1a4.port_a_logical_ram_width = 32;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.ram_block_type = "auto";
defparam ram_block1a4.mem_init0 = "79E89849B2238B9BB6E73FE43D9BC8C166A1F9C0F6BA1EAA08CF4554B8D8634A";

cyclonev_ram_block ram_block1a12(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a12_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a12.clk0_core_clock_enable = "ena0";
defparam ram_block1a12.clk0_input_clock_enable = "ena0";
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.init_file = "processor_cpu_ociram_default_contents.mif";
defparam ram_block1a12.init_file_layout = "port_a";
defparam ram_block1a12.logical_ram_name = "processor_cpu:cpu|processor_cpu_nios2_oci:the_processor_cpu_nios2_oci|processor_cpu_nios2_ocimem:the_processor_cpu_nios2_ocimem|processor_cpu_ociram_sp_ram_module:processor_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_4qe1:auto_generated|ALTSYNCRAM";
defparam ram_block1a12.operation_mode = "single_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 8;
defparam ram_block1a12.port_a_byte_enable_mask_width = 1;
defparam ram_block1a12.port_a_byte_size = 1;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 255;
defparam ram_block1a12.port_a_logical_ram_depth = 256;
defparam ram_block1a12.port_a_logical_ram_width = 32;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a12.ram_block_type = "auto";
defparam ram_block1a12.mem_init0 = "CAFE8146F9752B2065A8CED2B02561410CA1B76131DB11AC039226CDD69946D0";

cyclonev_ram_block ram_block1a28(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[28]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a28_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a28.clk0_core_clock_enable = "ena0";
defparam ram_block1a28.clk0_input_clock_enable = "ena0";
defparam ram_block1a28.data_interleave_offset_in_bits = 1;
defparam ram_block1a28.data_interleave_width_in_bits = 1;
defparam ram_block1a28.init_file = "processor_cpu_ociram_default_contents.mif";
defparam ram_block1a28.init_file_layout = "port_a";
defparam ram_block1a28.logical_ram_name = "processor_cpu:cpu|processor_cpu_nios2_oci:the_processor_cpu_nios2_oci|processor_cpu_nios2_ocimem:the_processor_cpu_nios2_ocimem|processor_cpu_ociram_sp_ram_module:processor_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_4qe1:auto_generated|ALTSYNCRAM";
defparam ram_block1a28.operation_mode = "single_port";
defparam ram_block1a28.port_a_address_clear = "none";
defparam ram_block1a28.port_a_address_width = 8;
defparam ram_block1a28.port_a_byte_enable_mask_width = 1;
defparam ram_block1a28.port_a_byte_size = 1;
defparam ram_block1a28.port_a_data_out_clear = "none";
defparam ram_block1a28.port_a_data_out_clock = "none";
defparam ram_block1a28.port_a_data_width = 1;
defparam ram_block1a28.port_a_first_address = 0;
defparam ram_block1a28.port_a_first_bit_number = 28;
defparam ram_block1a28.port_a_last_address = 255;
defparam ram_block1a28.port_a_logical_ram_depth = 256;
defparam ram_block1a28.port_a_logical_ram_width = 32;
defparam ram_block1a28.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a28.ram_block_type = "auto";
defparam ram_block1a28.mem_init0 = "A2230993CF91AB682BECD42F86F5803561257952176173A74D3B1FCD6A1E419D";

cyclonev_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a6_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a6.clk0_core_clock_enable = "ena0";
defparam ram_block1a6.clk0_input_clock_enable = "ena0";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.init_file = "processor_cpu_ociram_default_contents.mif";
defparam ram_block1a6.init_file_layout = "port_a";
defparam ram_block1a6.logical_ram_name = "processor_cpu:cpu|processor_cpu_nios2_oci:the_processor_cpu_nios2_oci|processor_cpu_nios2_ocimem:the_processor_cpu_nios2_ocimem|processor_cpu_ociram_sp_ram_module:processor_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_4qe1:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.operation_mode = "single_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 8;
defparam ram_block1a6.port_a_byte_enable_mask_width = 1;
defparam ram_block1a6.port_a_byte_size = 1;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 255;
defparam ram_block1a6.port_a_logical_ram_depth = 256;
defparam ram_block1a6.port_a_logical_ram_width = 32;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.ram_block_type = "auto";
defparam ram_block1a6.mem_init0 = "D88C8AC651B0172375610EAA646E019096C91D55B564B1D3FF42D916C0EE3F32";

cyclonev_ram_block ram_block1a22(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[22]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a22_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a22.clk0_core_clock_enable = "ena0";
defparam ram_block1a22.clk0_input_clock_enable = "ena0";
defparam ram_block1a22.data_interleave_offset_in_bits = 1;
defparam ram_block1a22.data_interleave_width_in_bits = 1;
defparam ram_block1a22.init_file = "processor_cpu_ociram_default_contents.mif";
defparam ram_block1a22.init_file_layout = "port_a";
defparam ram_block1a22.logical_ram_name = "processor_cpu:cpu|processor_cpu_nios2_oci:the_processor_cpu_nios2_oci|processor_cpu_nios2_ocimem:the_processor_cpu_nios2_ocimem|processor_cpu_ociram_sp_ram_module:processor_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_4qe1:auto_generated|ALTSYNCRAM";
defparam ram_block1a22.operation_mode = "single_port";
defparam ram_block1a22.port_a_address_clear = "none";
defparam ram_block1a22.port_a_address_width = 8;
defparam ram_block1a22.port_a_byte_enable_mask_width = 1;
defparam ram_block1a22.port_a_byte_size = 1;
defparam ram_block1a22.port_a_data_out_clear = "none";
defparam ram_block1a22.port_a_data_out_clock = "none";
defparam ram_block1a22.port_a_data_width = 1;
defparam ram_block1a22.port_a_first_address = 0;
defparam ram_block1a22.port_a_first_bit_number = 22;
defparam ram_block1a22.port_a_last_address = 255;
defparam ram_block1a22.port_a_logical_ram_depth = 256;
defparam ram_block1a22.port_a_logical_ram_width = 32;
defparam ram_block1a22.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a22.ram_block_type = "auto";
defparam ram_block1a22.mem_init0 = "A3D3B17971E078A0354875B91E2AA9D03DE4032006CE868643679723E8A2BD71";

cyclonev_ram_block ram_block1a14(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a14_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a14.clk0_core_clock_enable = "ena0";
defparam ram_block1a14.clk0_input_clock_enable = "ena0";
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.init_file = "processor_cpu_ociram_default_contents.mif";
defparam ram_block1a14.init_file_layout = "port_a";
defparam ram_block1a14.logical_ram_name = "processor_cpu:cpu|processor_cpu_nios2_oci:the_processor_cpu_nios2_oci|processor_cpu_nios2_ocimem:the_processor_cpu_nios2_ocimem|processor_cpu_ociram_sp_ram_module:processor_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_4qe1:auto_generated|ALTSYNCRAM";
defparam ram_block1a14.operation_mode = "single_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 8;
defparam ram_block1a14.port_a_byte_enable_mask_width = 1;
defparam ram_block1a14.port_a_byte_size = 1;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 255;
defparam ram_block1a14.port_a_logical_ram_depth = 256;
defparam ram_block1a14.port_a_logical_ram_width = 32;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a14.ram_block_type = "auto";
defparam ram_block1a14.mem_init0 = "3E15CCDE46521E7FCEBD107E14CF06B37D5ED68D563B69BD6DFD933781FE4DAE";

cyclonev_ram_block ram_block1a30(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[30]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a30_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a30.clk0_core_clock_enable = "ena0";
defparam ram_block1a30.clk0_input_clock_enable = "ena0";
defparam ram_block1a30.data_interleave_offset_in_bits = 1;
defparam ram_block1a30.data_interleave_width_in_bits = 1;
defparam ram_block1a30.init_file = "processor_cpu_ociram_default_contents.mif";
defparam ram_block1a30.init_file_layout = "port_a";
defparam ram_block1a30.logical_ram_name = "processor_cpu:cpu|processor_cpu_nios2_oci:the_processor_cpu_nios2_oci|processor_cpu_nios2_ocimem:the_processor_cpu_nios2_ocimem|processor_cpu_ociram_sp_ram_module:processor_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_4qe1:auto_generated|ALTSYNCRAM";
defparam ram_block1a30.operation_mode = "single_port";
defparam ram_block1a30.port_a_address_clear = "none";
defparam ram_block1a30.port_a_address_width = 8;
defparam ram_block1a30.port_a_byte_enable_mask_width = 1;
defparam ram_block1a30.port_a_byte_size = 1;
defparam ram_block1a30.port_a_data_out_clear = "none";
defparam ram_block1a30.port_a_data_out_clock = "none";
defparam ram_block1a30.port_a_data_width = 1;
defparam ram_block1a30.port_a_first_address = 0;
defparam ram_block1a30.port_a_first_bit_number = 30;
defparam ram_block1a30.port_a_last_address = 255;
defparam ram_block1a30.port_a_logical_ram_depth = 256;
defparam ram_block1a30.port_a_logical_ram_width = 32;
defparam ram_block1a30.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a30.ram_block_type = "auto";
defparam ram_block1a30.mem_init0 = "0D1DCE468A1830B27E519D02FAF7E48644C58296B6B82905784832211BF786B3";

cyclonev_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a7_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a7.clk0_core_clock_enable = "ena0";
defparam ram_block1a7.clk0_input_clock_enable = "ena0";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.init_file = "processor_cpu_ociram_default_contents.mif";
defparam ram_block1a7.init_file_layout = "port_a";
defparam ram_block1a7.logical_ram_name = "processor_cpu:cpu|processor_cpu_nios2_oci:the_processor_cpu_nios2_oci|processor_cpu_nios2_ocimem:the_processor_cpu_nios2_ocimem|processor_cpu_ociram_sp_ram_module:processor_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_4qe1:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.operation_mode = "single_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 8;
defparam ram_block1a7.port_a_byte_enable_mask_width = 1;
defparam ram_block1a7.port_a_byte_size = 1;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 255;
defparam ram_block1a7.port_a_logical_ram_depth = 256;
defparam ram_block1a7.port_a_logical_ram_width = 32;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.ram_block_type = "auto";
defparam ram_block1a7.mem_init0 = "809042A238CD1915199CC77B204E9890128E2108FD03AF3CD2C8AA6D944402B8";

cyclonev_ram_block ram_block1a23(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[23]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a23_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a23.clk0_core_clock_enable = "ena0";
defparam ram_block1a23.clk0_input_clock_enable = "ena0";
defparam ram_block1a23.data_interleave_offset_in_bits = 1;
defparam ram_block1a23.data_interleave_width_in_bits = 1;
defparam ram_block1a23.init_file = "processor_cpu_ociram_default_contents.mif";
defparam ram_block1a23.init_file_layout = "port_a";
defparam ram_block1a23.logical_ram_name = "processor_cpu:cpu|processor_cpu_nios2_oci:the_processor_cpu_nios2_oci|processor_cpu_nios2_ocimem:the_processor_cpu_nios2_ocimem|processor_cpu_ociram_sp_ram_module:processor_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_4qe1:auto_generated|ALTSYNCRAM";
defparam ram_block1a23.operation_mode = "single_port";
defparam ram_block1a23.port_a_address_clear = "none";
defparam ram_block1a23.port_a_address_width = 8;
defparam ram_block1a23.port_a_byte_enable_mask_width = 1;
defparam ram_block1a23.port_a_byte_size = 1;
defparam ram_block1a23.port_a_data_out_clear = "none";
defparam ram_block1a23.port_a_data_out_clock = "none";
defparam ram_block1a23.port_a_data_width = 1;
defparam ram_block1a23.port_a_first_address = 0;
defparam ram_block1a23.port_a_first_bit_number = 23;
defparam ram_block1a23.port_a_last_address = 255;
defparam ram_block1a23.port_a_logical_ram_depth = 256;
defparam ram_block1a23.port_a_logical_ram_width = 32;
defparam ram_block1a23.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a23.ram_block_type = "auto";
defparam ram_block1a23.mem_init0 = "F2FF32884A75FB4E414BCC5ED0D90F02E051607E458649819209FE2B47FD2FEC";

cyclonev_ram_block ram_block1a15(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a15_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a15.clk0_core_clock_enable = "ena0";
defparam ram_block1a15.clk0_input_clock_enable = "ena0";
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.init_file = "processor_cpu_ociram_default_contents.mif";
defparam ram_block1a15.init_file_layout = "port_a";
defparam ram_block1a15.logical_ram_name = "processor_cpu:cpu|processor_cpu_nios2_oci:the_processor_cpu_nios2_oci|processor_cpu_nios2_ocimem:the_processor_cpu_nios2_ocimem|processor_cpu_ociram_sp_ram_module:processor_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_4qe1:auto_generated|ALTSYNCRAM";
defparam ram_block1a15.operation_mode = "single_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 8;
defparam ram_block1a15.port_a_byte_enable_mask_width = 1;
defparam ram_block1a15.port_a_byte_size = 1;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 255;
defparam ram_block1a15.port_a_logical_ram_depth = 256;
defparam ram_block1a15.port_a_logical_ram_width = 32;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a15.ram_block_type = "auto";
defparam ram_block1a15.mem_init0 = "E454C43F0A08EDEA0EE78B116A19AFE6DB876AD24EC242817DED2798F34B1778";

cyclonev_ram_block ram_block1a31(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[31]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a31_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a31.clk0_core_clock_enable = "ena0";
defparam ram_block1a31.clk0_input_clock_enable = "ena0";
defparam ram_block1a31.data_interleave_offset_in_bits = 1;
defparam ram_block1a31.data_interleave_width_in_bits = 1;
defparam ram_block1a31.init_file = "processor_cpu_ociram_default_contents.mif";
defparam ram_block1a31.init_file_layout = "port_a";
defparam ram_block1a31.logical_ram_name = "processor_cpu:cpu|processor_cpu_nios2_oci:the_processor_cpu_nios2_oci|processor_cpu_nios2_ocimem:the_processor_cpu_nios2_ocimem|processor_cpu_ociram_sp_ram_module:processor_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_4qe1:auto_generated|ALTSYNCRAM";
defparam ram_block1a31.operation_mode = "single_port";
defparam ram_block1a31.port_a_address_clear = "none";
defparam ram_block1a31.port_a_address_width = 8;
defparam ram_block1a31.port_a_byte_enable_mask_width = 1;
defparam ram_block1a31.port_a_byte_size = 1;
defparam ram_block1a31.port_a_data_out_clear = "none";
defparam ram_block1a31.port_a_data_out_clock = "none";
defparam ram_block1a31.port_a_data_width = 1;
defparam ram_block1a31.port_a_first_address = 0;
defparam ram_block1a31.port_a_first_bit_number = 31;
defparam ram_block1a31.port_a_last_address = 255;
defparam ram_block1a31.port_a_logical_ram_depth = 256;
defparam ram_block1a31.port_a_logical_ram_width = 32;
defparam ram_block1a31.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a31.ram_block_type = "auto";
defparam ram_block1a31.mem_init0 = "8C39BEA8FC3C6D2B053FC6729A29ACA3A834D004F11037B3A1BC2994A7C386B6";

cyclonev_ram_block ram_block1a11(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a11_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a11.clk0_core_clock_enable = "ena0";
defparam ram_block1a11.clk0_input_clock_enable = "ena0";
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.init_file = "processor_cpu_ociram_default_contents.mif";
defparam ram_block1a11.init_file_layout = "port_a";
defparam ram_block1a11.logical_ram_name = "processor_cpu:cpu|processor_cpu_nios2_oci:the_processor_cpu_nios2_oci|processor_cpu_nios2_ocimem:the_processor_cpu_nios2_ocimem|processor_cpu_ociram_sp_ram_module:processor_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_4qe1:auto_generated|ALTSYNCRAM";
defparam ram_block1a11.operation_mode = "single_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 8;
defparam ram_block1a11.port_a_byte_enable_mask_width = 1;
defparam ram_block1a11.port_a_byte_size = 1;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 255;
defparam ram_block1a11.port_a_logical_ram_depth = 256;
defparam ram_block1a11.port_a_logical_ram_width = 32;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a11.ram_block_type = "auto";
defparam ram_block1a11.mem_init0 = "88E515FCA96491A7760B8047458582F91DAF2659A83C0CB059FF298547328EDE";

cyclonev_ram_block ram_block1a27(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[27]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a27_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a27.clk0_core_clock_enable = "ena0";
defparam ram_block1a27.clk0_input_clock_enable = "ena0";
defparam ram_block1a27.data_interleave_offset_in_bits = 1;
defparam ram_block1a27.data_interleave_width_in_bits = 1;
defparam ram_block1a27.init_file = "processor_cpu_ociram_default_contents.mif";
defparam ram_block1a27.init_file_layout = "port_a";
defparam ram_block1a27.logical_ram_name = "processor_cpu:cpu|processor_cpu_nios2_oci:the_processor_cpu_nios2_oci|processor_cpu_nios2_ocimem:the_processor_cpu_nios2_ocimem|processor_cpu_ociram_sp_ram_module:processor_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_4qe1:auto_generated|ALTSYNCRAM";
defparam ram_block1a27.operation_mode = "single_port";
defparam ram_block1a27.port_a_address_clear = "none";
defparam ram_block1a27.port_a_address_width = 8;
defparam ram_block1a27.port_a_byte_enable_mask_width = 1;
defparam ram_block1a27.port_a_byte_size = 1;
defparam ram_block1a27.port_a_data_out_clear = "none";
defparam ram_block1a27.port_a_data_out_clock = "none";
defparam ram_block1a27.port_a_data_width = 1;
defparam ram_block1a27.port_a_first_address = 0;
defparam ram_block1a27.port_a_first_bit_number = 27;
defparam ram_block1a27.port_a_last_address = 255;
defparam ram_block1a27.port_a_logical_ram_depth = 256;
defparam ram_block1a27.port_a_logical_ram_width = 32;
defparam ram_block1a27.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a27.ram_block_type = "auto";
defparam ram_block1a27.mem_init0 = "FB552A1D483607D3E50925BCD213C99CC386063369FA8A9CCF970F9F9D9061D7";

cyclonev_ram_block ram_block1a10(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a10_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a10.clk0_core_clock_enable = "ena0";
defparam ram_block1a10.clk0_input_clock_enable = "ena0";
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.init_file = "processor_cpu_ociram_default_contents.mif";
defparam ram_block1a10.init_file_layout = "port_a";
defparam ram_block1a10.logical_ram_name = "processor_cpu:cpu|processor_cpu_nios2_oci:the_processor_cpu_nios2_oci|processor_cpu_nios2_ocimem:the_processor_cpu_nios2_ocimem|processor_cpu_ociram_sp_ram_module:processor_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_4qe1:auto_generated|ALTSYNCRAM";
defparam ram_block1a10.operation_mode = "single_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 8;
defparam ram_block1a10.port_a_byte_enable_mask_width = 1;
defparam ram_block1a10.port_a_byte_size = 1;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 255;
defparam ram_block1a10.port_a_logical_ram_depth = 256;
defparam ram_block1a10.port_a_logical_ram_width = 32;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a10.ram_block_type = "auto";
defparam ram_block1a10.mem_init0 = "87C0D5782816FE7CE5847E0EC072EE77BF6263BECDFF886CA05DEE9D9BCB0525";

cyclonev_ram_block ram_block1a26(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[26]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a26_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a26.clk0_core_clock_enable = "ena0";
defparam ram_block1a26.clk0_input_clock_enable = "ena0";
defparam ram_block1a26.data_interleave_offset_in_bits = 1;
defparam ram_block1a26.data_interleave_width_in_bits = 1;
defparam ram_block1a26.init_file = "processor_cpu_ociram_default_contents.mif";
defparam ram_block1a26.init_file_layout = "port_a";
defparam ram_block1a26.logical_ram_name = "processor_cpu:cpu|processor_cpu_nios2_oci:the_processor_cpu_nios2_oci|processor_cpu_nios2_ocimem:the_processor_cpu_nios2_ocimem|processor_cpu_ociram_sp_ram_module:processor_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_4qe1:auto_generated|ALTSYNCRAM";
defparam ram_block1a26.operation_mode = "single_port";
defparam ram_block1a26.port_a_address_clear = "none";
defparam ram_block1a26.port_a_address_width = 8;
defparam ram_block1a26.port_a_byte_enable_mask_width = 1;
defparam ram_block1a26.port_a_byte_size = 1;
defparam ram_block1a26.port_a_data_out_clear = "none";
defparam ram_block1a26.port_a_data_out_clock = "none";
defparam ram_block1a26.port_a_data_width = 1;
defparam ram_block1a26.port_a_first_address = 0;
defparam ram_block1a26.port_a_first_bit_number = 26;
defparam ram_block1a26.port_a_last_address = 255;
defparam ram_block1a26.port_a_logical_ram_depth = 256;
defparam ram_block1a26.port_a_logical_ram_width = 32;
defparam ram_block1a26.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a26.ram_block_type = "auto";
defparam ram_block1a26.mem_init0 = "2B4C4C58C3FB8AF5BED936D1221A104CAA70AAD5276393433DE7BD3DB21479F9";

cyclonev_ram_block ram_block1a25(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[25]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a25_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a25.clk0_core_clock_enable = "ena0";
defparam ram_block1a25.clk0_input_clock_enable = "ena0";
defparam ram_block1a25.data_interleave_offset_in_bits = 1;
defparam ram_block1a25.data_interleave_width_in_bits = 1;
defparam ram_block1a25.init_file = "processor_cpu_ociram_default_contents.mif";
defparam ram_block1a25.init_file_layout = "port_a";
defparam ram_block1a25.logical_ram_name = "processor_cpu:cpu|processor_cpu_nios2_oci:the_processor_cpu_nios2_oci|processor_cpu_nios2_ocimem:the_processor_cpu_nios2_ocimem|processor_cpu_ociram_sp_ram_module:processor_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_4qe1:auto_generated|ALTSYNCRAM";
defparam ram_block1a25.operation_mode = "single_port";
defparam ram_block1a25.port_a_address_clear = "none";
defparam ram_block1a25.port_a_address_width = 8;
defparam ram_block1a25.port_a_byte_enable_mask_width = 1;
defparam ram_block1a25.port_a_byte_size = 1;
defparam ram_block1a25.port_a_data_out_clear = "none";
defparam ram_block1a25.port_a_data_out_clock = "none";
defparam ram_block1a25.port_a_data_width = 1;
defparam ram_block1a25.port_a_first_address = 0;
defparam ram_block1a25.port_a_first_bit_number = 25;
defparam ram_block1a25.port_a_last_address = 255;
defparam ram_block1a25.port_a_logical_ram_depth = 256;
defparam ram_block1a25.port_a_logical_ram_width = 32;
defparam ram_block1a25.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a25.ram_block_type = "auto";
defparam ram_block1a25.mem_init0 = "87894BF09AAB5618DC7D301FAFF1AB6CCC1AFF1791A2DF6D87C73D4D19C5D4FC";

cyclonev_ram_block ram_block1a9(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a9_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a9.clk0_core_clock_enable = "ena0";
defparam ram_block1a9.clk0_input_clock_enable = "ena0";
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.init_file = "processor_cpu_ociram_default_contents.mif";
defparam ram_block1a9.init_file_layout = "port_a";
defparam ram_block1a9.logical_ram_name = "processor_cpu:cpu|processor_cpu_nios2_oci:the_processor_cpu_nios2_oci|processor_cpu_nios2_ocimem:the_processor_cpu_nios2_ocimem|processor_cpu_ociram_sp_ram_module:processor_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_4qe1:auto_generated|ALTSYNCRAM";
defparam ram_block1a9.operation_mode = "single_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 8;
defparam ram_block1a9.port_a_byte_enable_mask_width = 1;
defparam ram_block1a9.port_a_byte_size = 1;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 255;
defparam ram_block1a9.port_a_logical_ram_depth = 256;
defparam ram_block1a9.port_a_logical_ram_width = 32;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a9.ram_block_type = "auto";
defparam ram_block1a9.mem_init0 = "8612C41166A7972AFBFFC4A72AA1DEC34D8048511E87B0B1E74FD4F920180336";

cyclonev_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a3_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a3.clk0_core_clock_enable = "ena0";
defparam ram_block1a3.clk0_input_clock_enable = "ena0";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.init_file = "processor_cpu_ociram_default_contents.mif";
defparam ram_block1a3.init_file_layout = "port_a";
defparam ram_block1a3.logical_ram_name = "processor_cpu:cpu|processor_cpu_nios2_oci:the_processor_cpu_nios2_oci|processor_cpu_nios2_ocimem:the_processor_cpu_nios2_ocimem|processor_cpu_ociram_sp_ram_module:processor_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_4qe1:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.operation_mode = "single_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 8;
defparam ram_block1a3.port_a_byte_enable_mask_width = 1;
defparam ram_block1a3.port_a_byte_size = 1;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 255;
defparam ram_block1a3.port_a_logical_ram_depth = 256;
defparam ram_block1a3.port_a_logical_ram_width = 32;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.ram_block_type = "auto";
defparam ram_block1a3.mem_init0 = "E633C4C82AD564200DDC93F4E4FCFE0F10D3E8843064AB49598E95C35A062282";

cyclonev_ram_block ram_block1a18(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[18]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a18_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a18.clk0_core_clock_enable = "ena0";
defparam ram_block1a18.clk0_input_clock_enable = "ena0";
defparam ram_block1a18.data_interleave_offset_in_bits = 1;
defparam ram_block1a18.data_interleave_width_in_bits = 1;
defparam ram_block1a18.init_file = "processor_cpu_ociram_default_contents.mif";
defparam ram_block1a18.init_file_layout = "port_a";
defparam ram_block1a18.logical_ram_name = "processor_cpu:cpu|processor_cpu_nios2_oci:the_processor_cpu_nios2_oci|processor_cpu_nios2_ocimem:the_processor_cpu_nios2_ocimem|processor_cpu_ociram_sp_ram_module:processor_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_4qe1:auto_generated|ALTSYNCRAM";
defparam ram_block1a18.operation_mode = "single_port";
defparam ram_block1a18.port_a_address_clear = "none";
defparam ram_block1a18.port_a_address_width = 8;
defparam ram_block1a18.port_a_byte_enable_mask_width = 1;
defparam ram_block1a18.port_a_byte_size = 1;
defparam ram_block1a18.port_a_data_out_clear = "none";
defparam ram_block1a18.port_a_data_out_clock = "none";
defparam ram_block1a18.port_a_data_width = 1;
defparam ram_block1a18.port_a_first_address = 0;
defparam ram_block1a18.port_a_first_bit_number = 18;
defparam ram_block1a18.port_a_last_address = 255;
defparam ram_block1a18.port_a_logical_ram_depth = 256;
defparam ram_block1a18.port_a_logical_ram_width = 32;
defparam ram_block1a18.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a18.ram_block_type = "auto";
defparam ram_block1a18.mem_init0 = "DEF2B79C2B0A6D738AD7EB2EFDC138C31CA5C1478DB6AE9DF5012164CC68E510";

cyclonev_ram_block ram_block1a17(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[17]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a17_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a17.clk0_core_clock_enable = "ena0";
defparam ram_block1a17.clk0_input_clock_enable = "ena0";
defparam ram_block1a17.data_interleave_offset_in_bits = 1;
defparam ram_block1a17.data_interleave_width_in_bits = 1;
defparam ram_block1a17.init_file = "processor_cpu_ociram_default_contents.mif";
defparam ram_block1a17.init_file_layout = "port_a";
defparam ram_block1a17.logical_ram_name = "processor_cpu:cpu|processor_cpu_nios2_oci:the_processor_cpu_nios2_oci|processor_cpu_nios2_ocimem:the_processor_cpu_nios2_ocimem|processor_cpu_ociram_sp_ram_module:processor_cpu_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_4qe1:auto_generated|ALTSYNCRAM";
defparam ram_block1a17.operation_mode = "single_port";
defparam ram_block1a17.port_a_address_clear = "none";
defparam ram_block1a17.port_a_address_width = 8;
defparam ram_block1a17.port_a_byte_enable_mask_width = 1;
defparam ram_block1a17.port_a_byte_size = 1;
defparam ram_block1a17.port_a_data_out_clear = "none";
defparam ram_block1a17.port_a_data_out_clock = "none";
defparam ram_block1a17.port_a_data_width = 1;
defparam ram_block1a17.port_a_first_address = 0;
defparam ram_block1a17.port_a_first_bit_number = 17;
defparam ram_block1a17.port_a_last_address = 255;
defparam ram_block1a17.port_a_logical_ram_depth = 256;
defparam ram_block1a17.port_a_logical_ram_width = 32;
defparam ram_block1a17.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a17.ram_block_type = "auto";
defparam ram_block1a17.mem_init0 = "C1F7B73EE93A06E9824DC9DAEC9FDFADDB2ACDCFC8DEFA542138FA129ED25A18";

endmodule

module processor_processor_cpu_register_bank_a_module (
	q_b_5,
	q_b_4,
	q_b_6,
	q_b_16,
	q_b_15,
	q_b_14,
	q_b_13,
	q_b_12,
	q_b_11,
	q_b_10,
	q_b_9,
	q_b_8,
	q_b_7,
	q_b_3,
	q_b_2,
	q_b_0,
	q_b_29,
	q_b_27,
	q_b_28,
	q_b_30,
	q_b_31,
	q_b_1,
	q_b_311,
	q_b_17,
	q_b_301,
	q_b_18,
	q_b_291,
	q_b_19,
	q_b_281,
	q_b_24,
	q_b_21,
	q_b_20,
	q_b_22,
	q_b_23,
	q_b_271,
	q_b_26,
	q_b_25,
	W_stall,
	M_wr_data_unfiltered_5,
	M_wr_data_unfiltered_15,
	M_wr_data_unfiltered_14,
	M_wr_data_unfiltered_13,
	M_wr_data_unfiltered_12,
	M_wr_data_unfiltered_11,
	M_wr_data_unfiltered_9,
	M_wr_data_unfiltered_7,
	M_wr_data_unfiltered_3,
	M_wr_data_unfiltered_1,
	M_wr_data_unfiltered_0,
	M_dst_regnum_4,
	M_wr_dst_reg,
	M_dst_regnum_0,
	M_dst_regnum_1,
	M_dst_regnum_2,
	M_dst_regnum_3,
	M_wr_data_unfiltered_4,
	M_wr_data_unfiltered_6,
	M_wr_data_unfiltered_16,
	M_wr_data_unfiltered_10,
	M_wr_data_unfiltered_8,
	M_wr_data_unfiltered_2,
	M_wr_data_unfiltered_31,
	M_wr_data_unfiltered_17,
	M_wr_data_unfiltered_30,
	M_wr_data_unfiltered_29,
	M_wr_data_unfiltered_21,
	M_wr_data_unfiltered_19,
	M_wr_data_unfiltered_18,
	M_wr_data_unfiltered_23,
	M_wr_data_unfiltered_27,
	M_wr_data_unfiltered_25,
	M_wr_data_unfiltered_24,
	M_wr_data_unfiltered_20,
	M_wr_data_unfiltered_28,
	M_wr_data_unfiltered_22,
	M_wr_data_unfiltered_26,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_5;
output 	q_b_4;
output 	q_b_6;
output 	q_b_16;
output 	q_b_15;
output 	q_b_14;
output 	q_b_13;
output 	q_b_12;
output 	q_b_11;
output 	q_b_10;
output 	q_b_9;
output 	q_b_8;
output 	q_b_7;
output 	q_b_3;
output 	q_b_2;
output 	q_b_0;
input 	q_b_29;
input 	q_b_27;
input 	q_b_28;
input 	q_b_30;
input 	q_b_31;
output 	q_b_1;
output 	q_b_311;
output 	q_b_17;
output 	q_b_301;
output 	q_b_18;
output 	q_b_291;
output 	q_b_19;
output 	q_b_281;
output 	q_b_24;
output 	q_b_21;
output 	q_b_20;
output 	q_b_22;
output 	q_b_23;
output 	q_b_271;
output 	q_b_26;
output 	q_b_25;
input 	W_stall;
input 	M_wr_data_unfiltered_5;
input 	M_wr_data_unfiltered_15;
input 	M_wr_data_unfiltered_14;
input 	M_wr_data_unfiltered_13;
input 	M_wr_data_unfiltered_12;
input 	M_wr_data_unfiltered_11;
input 	M_wr_data_unfiltered_9;
input 	M_wr_data_unfiltered_7;
input 	M_wr_data_unfiltered_3;
input 	M_wr_data_unfiltered_1;
input 	M_wr_data_unfiltered_0;
input 	M_dst_regnum_4;
input 	M_wr_dst_reg;
input 	M_dst_regnum_0;
input 	M_dst_regnum_1;
input 	M_dst_regnum_2;
input 	M_dst_regnum_3;
input 	M_wr_data_unfiltered_4;
input 	M_wr_data_unfiltered_6;
input 	M_wr_data_unfiltered_16;
input 	M_wr_data_unfiltered_10;
input 	M_wr_data_unfiltered_8;
input 	M_wr_data_unfiltered_2;
input 	M_wr_data_unfiltered_31;
input 	M_wr_data_unfiltered_17;
input 	M_wr_data_unfiltered_30;
input 	M_wr_data_unfiltered_29;
input 	M_wr_data_unfiltered_21;
input 	M_wr_data_unfiltered_19;
input 	M_wr_data_unfiltered_18;
input 	M_wr_data_unfiltered_23;
input 	M_wr_data_unfiltered_27;
input 	M_wr_data_unfiltered_25;
input 	M_wr_data_unfiltered_24;
input 	M_wr_data_unfiltered_20;
input 	M_wr_data_unfiltered_28;
input 	M_wr_data_unfiltered_22;
input 	M_wr_data_unfiltered_26;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



processor_altsyncram_4 the_altsyncram(
	.q_b({q_b_311,q_b_301,q_b_291,q_b_281,q_b_271,q_b_26,q_b_25,q_b_24,q_b_23,q_b_22,q_b_21,q_b_20,q_b_19,q_b_18,q_b_17,q_b_16,q_b_15,q_b_14,q_b_13,q_b_12,q_b_11,q_b_10,q_b_9,q_b_8,q_b_7,q_b_6,q_b_5,q_b_4,q_b_3,q_b_2,q_b_1,q_b_0}),
	.address_b({gnd,gnd,gnd,gnd,q_b_31,q_b_30,q_b_29,q_b_28,q_b_27}),
	.rden_b(W_stall),
	.data_a({M_wr_data_unfiltered_31,M_wr_data_unfiltered_30,M_wr_data_unfiltered_29,M_wr_data_unfiltered_28,M_wr_data_unfiltered_27,M_wr_data_unfiltered_26,M_wr_data_unfiltered_25,M_wr_data_unfiltered_24,M_wr_data_unfiltered_23,M_wr_data_unfiltered_22,M_wr_data_unfiltered_21,
M_wr_data_unfiltered_20,M_wr_data_unfiltered_19,M_wr_data_unfiltered_18,M_wr_data_unfiltered_17,M_wr_data_unfiltered_16,M_wr_data_unfiltered_15,M_wr_data_unfiltered_14,M_wr_data_unfiltered_13,M_wr_data_unfiltered_12,M_wr_data_unfiltered_11,M_wr_data_unfiltered_10,
M_wr_data_unfiltered_9,M_wr_data_unfiltered_8,M_wr_data_unfiltered_7,M_wr_data_unfiltered_6,M_wr_data_unfiltered_5,M_wr_data_unfiltered_4,M_wr_data_unfiltered_3,M_wr_data_unfiltered_2,M_wr_data_unfiltered_1,M_wr_data_unfiltered_0}),
	.address_a({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,M_dst_regnum_4,M_dst_regnum_3,M_dst_regnum_2,M_dst_regnum_1,M_dst_regnum_0}),
	.wren_a(M_wr_dst_reg),
	.clock0(clk_clk));

endmodule

module processor_altsyncram_4 (
	q_b,
	address_b,
	rden_b,
	data_a,
	address_a,
	wren_a,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[31:0] q_b;
input 	[8:0] address_b;
input 	rden_b;
input 	[31:0] data_a;
input 	[12:0] address_a;
input 	wren_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



processor_altsyncram_44n1 auto_generated(
	.q_b({q_b[31],q_b[30],q_b[29],q_b[28],q_b[27],q_b[26],q_b[25],q_b[24],q_b[23],q_b[22],q_b[21],q_b[20],q_b[19],q_b[18],q_b[17],q_b[16],q_b[15],q_b[14],q_b[13],q_b[12],q_b[11],q_b[10],q_b[9],q_b[8],q_b[7],q_b[6],q_b[5],q_b[4],q_b[3],q_b[2],q_b[1],q_b[0]}),
	.address_b({address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.rden_b(rden_b),
	.data_a({data_a[31],data_a[30],data_a[29],data_a[28],data_a[27],data_a[26],data_a[25],data_a[24],data_a[23],data_a[22],data_a[21],data_a[20],data_a[19],data_a[18],data_a[17],data_a[16],data_a[15],data_a[14],data_a[13],data_a[12],data_a[11],data_a[10],data_a[9],data_a[8],data_a[7],data_a[6],data_a[5],data_a[4],data_a[3],data_a[2],data_a[1],data_a[0]}),
	.address_a({address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.wren_a(wren_a),
	.clock0(clock0));

endmodule

module processor_altsyncram_44n1 (
	q_b,
	address_b,
	rden_b,
	data_a,
	address_a,
	wren_a,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[31:0] q_b;
input 	[4:0] address_b;
input 	rden_b;
input 	[31:0] data_a;
input 	[4:0] address_a;
input 	wren_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a4_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a16_PORTBDATAOUT_bus;
wire [143:0] ram_block1a15_PORTBDATAOUT_bus;
wire [143:0] ram_block1a14_PORTBDATAOUT_bus;
wire [143:0] ram_block1a13_PORTBDATAOUT_bus;
wire [143:0] ram_block1a12_PORTBDATAOUT_bus;
wire [143:0] ram_block1a11_PORTBDATAOUT_bus;
wire [143:0] ram_block1a10_PORTBDATAOUT_bus;
wire [143:0] ram_block1a9_PORTBDATAOUT_bus;
wire [143:0] ram_block1a8_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;
wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a0_PORTBDATAOUT_bus;
wire [143:0] ram_block1a1_PORTBDATAOUT_bus;
wire [143:0] ram_block1a31_PORTBDATAOUT_bus;
wire [143:0] ram_block1a17_PORTBDATAOUT_bus;
wire [143:0] ram_block1a30_PORTBDATAOUT_bus;
wire [143:0] ram_block1a18_PORTBDATAOUT_bus;
wire [143:0] ram_block1a29_PORTBDATAOUT_bus;
wire [143:0] ram_block1a19_PORTBDATAOUT_bus;
wire [143:0] ram_block1a28_PORTBDATAOUT_bus;
wire [143:0] ram_block1a24_PORTBDATAOUT_bus;
wire [143:0] ram_block1a21_PORTBDATAOUT_bus;
wire [143:0] ram_block1a20_PORTBDATAOUT_bus;
wire [143:0] ram_block1a22_PORTBDATAOUT_bus;
wire [143:0] ram_block1a23_PORTBDATAOUT_bus;
wire [143:0] ram_block1a27_PORTBDATAOUT_bus;
wire [143:0] ram_block1a26_PORTBDATAOUT_bus;
wire [143:0] ram_block1a25_PORTBDATAOUT_bus;

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_b[16] = ram_block1a16_PORTBDATAOUT_bus[0];

assign q_b[15] = ram_block1a15_PORTBDATAOUT_bus[0];

assign q_b[14] = ram_block1a14_PORTBDATAOUT_bus[0];

assign q_b[13] = ram_block1a13_PORTBDATAOUT_bus[0];

assign q_b[12] = ram_block1a12_PORTBDATAOUT_bus[0];

assign q_b[11] = ram_block1a11_PORTBDATAOUT_bus[0];

assign q_b[10] = ram_block1a10_PORTBDATAOUT_bus[0];

assign q_b[9] = ram_block1a9_PORTBDATAOUT_bus[0];

assign q_b[8] = ram_block1a8_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_b[3] = ram_block1a3_PORTBDATAOUT_bus[0];

assign q_b[2] = ram_block1a2_PORTBDATAOUT_bus[0];

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

assign q_b[31] = ram_block1a31_PORTBDATAOUT_bus[0];

assign q_b[17] = ram_block1a17_PORTBDATAOUT_bus[0];

assign q_b[30] = ram_block1a30_PORTBDATAOUT_bus[0];

assign q_b[18] = ram_block1a18_PORTBDATAOUT_bus[0];

assign q_b[29] = ram_block1a29_PORTBDATAOUT_bus[0];

assign q_b[19] = ram_block1a19_PORTBDATAOUT_bus[0];

assign q_b[28] = ram_block1a28_PORTBDATAOUT_bus[0];

assign q_b[24] = ram_block1a24_PORTBDATAOUT_bus[0];

assign q_b[21] = ram_block1a21_PORTBDATAOUT_bus[0];

assign q_b[20] = ram_block1a20_PORTBDATAOUT_bus[0];

assign q_b[22] = ram_block1a22_PORTBDATAOUT_bus[0];

assign q_b[23] = ram_block1a23_PORTBDATAOUT_bus[0];

assign q_b[27] = ram_block1a27_PORTBDATAOUT_bus[0];

assign q_b[26] = ram_block1a26_PORTBDATAOUT_bus[0];

assign q_b[25] = ram_block1a25_PORTBDATAOUT_bus[0];

cyclonev_ram_block ram_block1a5(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.init_file = "processor_cpu_rf_ram_a.mif";
defparam ram_block1a5.init_file_layout = "port_b";
defparam ram_block1a5.logical_ram_name = "processor_cpu:cpu|processor_cpu_register_bank_a_module:processor_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_44n1:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "old";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 5;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 31;
defparam ram_block1a5.port_a_logical_ram_depth = 32;
defparam ram_block1a5.port_a_logical_ram_width = 32;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_address_clear = "none";
defparam ram_block1a5.port_b_address_clock = "clock0";
defparam ram_block1a5.port_b_address_width = 5;
defparam ram_block1a5.port_b_data_out_clear = "none";
defparam ram_block1a5.port_b_data_out_clock = "none";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 31;
defparam ram_block1a5.port_b_logical_ram_depth = 32;
defparam ram_block1a5.port_b_logical_ram_width = 32;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock0";
defparam ram_block1a5.ram_block_type = "auto";
defparam ram_block1a5.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a4(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.init_file = "processor_cpu_rf_ram_a.mif";
defparam ram_block1a4.init_file_layout = "port_b";
defparam ram_block1a4.logical_ram_name = "processor_cpu:cpu|processor_cpu_register_bank_a_module:processor_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_44n1:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "old";
defparam ram_block1a4.operation_mode = "dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 5;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 31;
defparam ram_block1a4.port_a_logical_ram_depth = 32;
defparam ram_block1a4.port_a_logical_ram_width = 32;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_address_clear = "none";
defparam ram_block1a4.port_b_address_clock = "clock0";
defparam ram_block1a4.port_b_address_width = 5;
defparam ram_block1a4.port_b_data_out_clear = "none";
defparam ram_block1a4.port_b_data_out_clock = "none";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 31;
defparam ram_block1a4.port_b_logical_ram_depth = 32;
defparam ram_block1a4.port_b_logical_ram_width = 32;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock0";
defparam ram_block1a4.ram_block_type = "auto";
defparam ram_block1a4.mem_init0 = "00000000";

cyclonev_ram_block ram_block1a6(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.init_file = "processor_cpu_rf_ram_a.mif";
defparam ram_block1a6.init_file_layout = "port_b";
defparam ram_block1a6.logical_ram_name = "processor_cpu:cpu|processor_cpu_register_bank_a_module:processor_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_44n1:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "old";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 5;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 31;
defparam ram_block1a6.port_a_logical_ram_depth = 32;
defparam ram_block1a6.port_a_logical_ram_width = 32;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_address_clear = "none";
defparam ram_block1a6.port_b_address_clock = "clock0";
defparam ram_block1a6.port_b_address_width = 5;
defparam ram_block1a6.port_b_data_out_clear = "none";
defparam ram_block1a6.port_b_data_out_clock = "none";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 31;
defparam ram_block1a6.port_b_logical_ram_depth = 32;
defparam ram_block1a6.port_b_logical_ram_width = 32;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock0";
defparam ram_block1a6.ram_block_type = "auto";
defparam ram_block1a6.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a16(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a16_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a16.data_interleave_offset_in_bits = 1;
defparam ram_block1a16.data_interleave_width_in_bits = 1;
defparam ram_block1a16.init_file = "processor_cpu_rf_ram_a.mif";
defparam ram_block1a16.init_file_layout = "port_b";
defparam ram_block1a16.logical_ram_name = "processor_cpu:cpu|processor_cpu_register_bank_a_module:processor_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_44n1:auto_generated|ALTSYNCRAM";
defparam ram_block1a16.mixed_port_feed_through_mode = "old";
defparam ram_block1a16.operation_mode = "dual_port";
defparam ram_block1a16.port_a_address_clear = "none";
defparam ram_block1a16.port_a_address_width = 5;
defparam ram_block1a16.port_a_data_out_clear = "none";
defparam ram_block1a16.port_a_data_out_clock = "none";
defparam ram_block1a16.port_a_data_width = 1;
defparam ram_block1a16.port_a_first_address = 0;
defparam ram_block1a16.port_a_first_bit_number = 16;
defparam ram_block1a16.port_a_last_address = 31;
defparam ram_block1a16.port_a_logical_ram_depth = 32;
defparam ram_block1a16.port_a_logical_ram_width = 32;
defparam ram_block1a16.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a16.port_b_address_clear = "none";
defparam ram_block1a16.port_b_address_clock = "clock0";
defparam ram_block1a16.port_b_address_width = 5;
defparam ram_block1a16.port_b_data_out_clear = "none";
defparam ram_block1a16.port_b_data_out_clock = "none";
defparam ram_block1a16.port_b_data_width = 1;
defparam ram_block1a16.port_b_first_address = 0;
defparam ram_block1a16.port_b_first_bit_number = 16;
defparam ram_block1a16.port_b_last_address = 31;
defparam ram_block1a16.port_b_logical_ram_depth = 32;
defparam ram_block1a16.port_b_logical_ram_width = 32;
defparam ram_block1a16.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a16.port_b_read_enable_clock = "clock0";
defparam ram_block1a16.ram_block_type = "auto";
defparam ram_block1a16.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a15(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a15_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.init_file = "processor_cpu_rf_ram_a.mif";
defparam ram_block1a15.init_file_layout = "port_b";
defparam ram_block1a15.logical_ram_name = "processor_cpu:cpu|processor_cpu_register_bank_a_module:processor_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_44n1:auto_generated|ALTSYNCRAM";
defparam ram_block1a15.mixed_port_feed_through_mode = "old";
defparam ram_block1a15.operation_mode = "dual_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 5;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 31;
defparam ram_block1a15.port_a_logical_ram_depth = 32;
defparam ram_block1a15.port_a_logical_ram_width = 32;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a15.port_b_address_clear = "none";
defparam ram_block1a15.port_b_address_clock = "clock0";
defparam ram_block1a15.port_b_address_width = 5;
defparam ram_block1a15.port_b_data_out_clear = "none";
defparam ram_block1a15.port_b_data_out_clock = "none";
defparam ram_block1a15.port_b_data_width = 1;
defparam ram_block1a15.port_b_first_address = 0;
defparam ram_block1a15.port_b_first_bit_number = 15;
defparam ram_block1a15.port_b_last_address = 31;
defparam ram_block1a15.port_b_logical_ram_depth = 32;
defparam ram_block1a15.port_b_logical_ram_width = 32;
defparam ram_block1a15.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a15.port_b_read_enable_clock = "clock0";
defparam ram_block1a15.ram_block_type = "auto";
defparam ram_block1a15.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a14(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a14_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.init_file = "processor_cpu_rf_ram_a.mif";
defparam ram_block1a14.init_file_layout = "port_b";
defparam ram_block1a14.logical_ram_name = "processor_cpu:cpu|processor_cpu_register_bank_a_module:processor_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_44n1:auto_generated|ALTSYNCRAM";
defparam ram_block1a14.mixed_port_feed_through_mode = "old";
defparam ram_block1a14.operation_mode = "dual_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 5;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 31;
defparam ram_block1a14.port_a_logical_ram_depth = 32;
defparam ram_block1a14.port_a_logical_ram_width = 32;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a14.port_b_address_clear = "none";
defparam ram_block1a14.port_b_address_clock = "clock0";
defparam ram_block1a14.port_b_address_width = 5;
defparam ram_block1a14.port_b_data_out_clear = "none";
defparam ram_block1a14.port_b_data_out_clock = "none";
defparam ram_block1a14.port_b_data_width = 1;
defparam ram_block1a14.port_b_first_address = 0;
defparam ram_block1a14.port_b_first_bit_number = 14;
defparam ram_block1a14.port_b_last_address = 31;
defparam ram_block1a14.port_b_logical_ram_depth = 32;
defparam ram_block1a14.port_b_logical_ram_width = 32;
defparam ram_block1a14.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a14.port_b_read_enable_clock = "clock0";
defparam ram_block1a14.ram_block_type = "auto";
defparam ram_block1a14.mem_init0 = "00000000";

cyclonev_ram_block ram_block1a13(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a13_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.init_file = "processor_cpu_rf_ram_a.mif";
defparam ram_block1a13.init_file_layout = "port_b";
defparam ram_block1a13.logical_ram_name = "processor_cpu:cpu|processor_cpu_register_bank_a_module:processor_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_44n1:auto_generated|ALTSYNCRAM";
defparam ram_block1a13.mixed_port_feed_through_mode = "old";
defparam ram_block1a13.operation_mode = "dual_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 5;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 31;
defparam ram_block1a13.port_a_logical_ram_depth = 32;
defparam ram_block1a13.port_a_logical_ram_width = 32;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a13.port_b_address_clear = "none";
defparam ram_block1a13.port_b_address_clock = "clock0";
defparam ram_block1a13.port_b_address_width = 5;
defparam ram_block1a13.port_b_data_out_clear = "none";
defparam ram_block1a13.port_b_data_out_clock = "none";
defparam ram_block1a13.port_b_data_width = 1;
defparam ram_block1a13.port_b_first_address = 0;
defparam ram_block1a13.port_b_first_bit_number = 13;
defparam ram_block1a13.port_b_last_address = 31;
defparam ram_block1a13.port_b_logical_ram_depth = 32;
defparam ram_block1a13.port_b_logical_ram_width = 32;
defparam ram_block1a13.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a13.port_b_read_enable_clock = "clock0";
defparam ram_block1a13.ram_block_type = "auto";
defparam ram_block1a13.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a12(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a12_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.init_file = "processor_cpu_rf_ram_a.mif";
defparam ram_block1a12.init_file_layout = "port_b";
defparam ram_block1a12.logical_ram_name = "processor_cpu:cpu|processor_cpu_register_bank_a_module:processor_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_44n1:auto_generated|ALTSYNCRAM";
defparam ram_block1a12.mixed_port_feed_through_mode = "old";
defparam ram_block1a12.operation_mode = "dual_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 5;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 31;
defparam ram_block1a12.port_a_logical_ram_depth = 32;
defparam ram_block1a12.port_a_logical_ram_width = 32;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a12.port_b_address_clear = "none";
defparam ram_block1a12.port_b_address_clock = "clock0";
defparam ram_block1a12.port_b_address_width = 5;
defparam ram_block1a12.port_b_data_out_clear = "none";
defparam ram_block1a12.port_b_data_out_clock = "none";
defparam ram_block1a12.port_b_data_width = 1;
defparam ram_block1a12.port_b_first_address = 0;
defparam ram_block1a12.port_b_first_bit_number = 12;
defparam ram_block1a12.port_b_last_address = 31;
defparam ram_block1a12.port_b_logical_ram_depth = 32;
defparam ram_block1a12.port_b_logical_ram_width = 32;
defparam ram_block1a12.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a12.port_b_read_enable_clock = "clock0";
defparam ram_block1a12.ram_block_type = "auto";
defparam ram_block1a12.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a11(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a11_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.init_file = "processor_cpu_rf_ram_a.mif";
defparam ram_block1a11.init_file_layout = "port_b";
defparam ram_block1a11.logical_ram_name = "processor_cpu:cpu|processor_cpu_register_bank_a_module:processor_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_44n1:auto_generated|ALTSYNCRAM";
defparam ram_block1a11.mixed_port_feed_through_mode = "old";
defparam ram_block1a11.operation_mode = "dual_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 5;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 31;
defparam ram_block1a11.port_a_logical_ram_depth = 32;
defparam ram_block1a11.port_a_logical_ram_width = 32;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a11.port_b_address_clear = "none";
defparam ram_block1a11.port_b_address_clock = "clock0";
defparam ram_block1a11.port_b_address_width = 5;
defparam ram_block1a11.port_b_data_out_clear = "none";
defparam ram_block1a11.port_b_data_out_clock = "none";
defparam ram_block1a11.port_b_data_width = 1;
defparam ram_block1a11.port_b_first_address = 0;
defparam ram_block1a11.port_b_first_bit_number = 11;
defparam ram_block1a11.port_b_last_address = 31;
defparam ram_block1a11.port_b_logical_ram_depth = 32;
defparam ram_block1a11.port_b_logical_ram_width = 32;
defparam ram_block1a11.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a11.port_b_read_enable_clock = "clock0";
defparam ram_block1a11.ram_block_type = "auto";
defparam ram_block1a11.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a10(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a10_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.init_file = "processor_cpu_rf_ram_a.mif";
defparam ram_block1a10.init_file_layout = "port_b";
defparam ram_block1a10.logical_ram_name = "processor_cpu:cpu|processor_cpu_register_bank_a_module:processor_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_44n1:auto_generated|ALTSYNCRAM";
defparam ram_block1a10.mixed_port_feed_through_mode = "old";
defparam ram_block1a10.operation_mode = "dual_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 5;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 31;
defparam ram_block1a10.port_a_logical_ram_depth = 32;
defparam ram_block1a10.port_a_logical_ram_width = 32;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a10.port_b_address_clear = "none";
defparam ram_block1a10.port_b_address_clock = "clock0";
defparam ram_block1a10.port_b_address_width = 5;
defparam ram_block1a10.port_b_data_out_clear = "none";
defparam ram_block1a10.port_b_data_out_clock = "none";
defparam ram_block1a10.port_b_data_width = 1;
defparam ram_block1a10.port_b_first_address = 0;
defparam ram_block1a10.port_b_first_bit_number = 10;
defparam ram_block1a10.port_b_last_address = 31;
defparam ram_block1a10.port_b_logical_ram_depth = 32;
defparam ram_block1a10.port_b_logical_ram_width = 32;
defparam ram_block1a10.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a10.port_b_read_enable_clock = "clock0";
defparam ram_block1a10.ram_block_type = "auto";
defparam ram_block1a10.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a9(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a9_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.init_file = "processor_cpu_rf_ram_a.mif";
defparam ram_block1a9.init_file_layout = "port_b";
defparam ram_block1a9.logical_ram_name = "processor_cpu:cpu|processor_cpu_register_bank_a_module:processor_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_44n1:auto_generated|ALTSYNCRAM";
defparam ram_block1a9.mixed_port_feed_through_mode = "old";
defparam ram_block1a9.operation_mode = "dual_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 5;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 31;
defparam ram_block1a9.port_a_logical_ram_depth = 32;
defparam ram_block1a9.port_a_logical_ram_width = 32;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a9.port_b_address_clear = "none";
defparam ram_block1a9.port_b_address_clock = "clock0";
defparam ram_block1a9.port_b_address_width = 5;
defparam ram_block1a9.port_b_data_out_clear = "none";
defparam ram_block1a9.port_b_data_out_clock = "none";
defparam ram_block1a9.port_b_data_width = 1;
defparam ram_block1a9.port_b_first_address = 0;
defparam ram_block1a9.port_b_first_bit_number = 9;
defparam ram_block1a9.port_b_last_address = 31;
defparam ram_block1a9.port_b_logical_ram_depth = 32;
defparam ram_block1a9.port_b_logical_ram_width = 32;
defparam ram_block1a9.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a9.port_b_read_enable_clock = "clock0";
defparam ram_block1a9.ram_block_type = "auto";
defparam ram_block1a9.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a8(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a8_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.init_file = "processor_cpu_rf_ram_a.mif";
defparam ram_block1a8.init_file_layout = "port_b";
defparam ram_block1a8.logical_ram_name = "processor_cpu:cpu|processor_cpu_register_bank_a_module:processor_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_44n1:auto_generated|ALTSYNCRAM";
defparam ram_block1a8.mixed_port_feed_through_mode = "old";
defparam ram_block1a8.operation_mode = "dual_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 5;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 31;
defparam ram_block1a8.port_a_logical_ram_depth = 32;
defparam ram_block1a8.port_a_logical_ram_width = 32;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a8.port_b_address_clear = "none";
defparam ram_block1a8.port_b_address_clock = "clock0";
defparam ram_block1a8.port_b_address_width = 5;
defparam ram_block1a8.port_b_data_out_clear = "none";
defparam ram_block1a8.port_b_data_out_clock = "none";
defparam ram_block1a8.port_b_data_width = 1;
defparam ram_block1a8.port_b_first_address = 0;
defparam ram_block1a8.port_b_first_bit_number = 8;
defparam ram_block1a8.port_b_last_address = 31;
defparam ram_block1a8.port_b_logical_ram_depth = 32;
defparam ram_block1a8.port_b_logical_ram_width = 32;
defparam ram_block1a8.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a8.port_b_read_enable_clock = "clock0";
defparam ram_block1a8.ram_block_type = "auto";
defparam ram_block1a8.mem_init0 = "00000000";

cyclonev_ram_block ram_block1a7(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.init_file = "processor_cpu_rf_ram_a.mif";
defparam ram_block1a7.init_file_layout = "port_b";
defparam ram_block1a7.logical_ram_name = "processor_cpu:cpu|processor_cpu_register_bank_a_module:processor_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_44n1:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "old";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 5;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 31;
defparam ram_block1a7.port_a_logical_ram_depth = 32;
defparam ram_block1a7.port_a_logical_ram_width = 32;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_address_clear = "none";
defparam ram_block1a7.port_b_address_clock = "clock0";
defparam ram_block1a7.port_b_address_width = 5;
defparam ram_block1a7.port_b_data_out_clear = "none";
defparam ram_block1a7.port_b_data_out_clock = "none";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 31;
defparam ram_block1a7.port_b_logical_ram_depth = 32;
defparam ram_block1a7.port_b_logical_ram_width = 32;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock0";
defparam ram_block1a7.ram_block_type = "auto";
defparam ram_block1a7.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a3(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.init_file = "processor_cpu_rf_ram_a.mif";
defparam ram_block1a3.init_file_layout = "port_b";
defparam ram_block1a3.logical_ram_name = "processor_cpu:cpu|processor_cpu_register_bank_a_module:processor_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_44n1:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "old";
defparam ram_block1a3.operation_mode = "dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 5;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 31;
defparam ram_block1a3.port_a_logical_ram_depth = 32;
defparam ram_block1a3.port_a_logical_ram_width = 32;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_address_clear = "none";
defparam ram_block1a3.port_b_address_clock = "clock0";
defparam ram_block1a3.port_b_address_width = 5;
defparam ram_block1a3.port_b_data_out_clear = "none";
defparam ram_block1a3.port_b_data_out_clock = "none";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 31;
defparam ram_block1a3.port_b_logical_ram_depth = 32;
defparam ram_block1a3.port_b_logical_ram_width = 32;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock0";
defparam ram_block1a3.ram_block_type = "auto";
defparam ram_block1a3.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a2(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.init_file = "processor_cpu_rf_ram_a.mif";
defparam ram_block1a2.init_file_layout = "port_b";
defparam ram_block1a2.logical_ram_name = "processor_cpu:cpu|processor_cpu_register_bank_a_module:processor_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_44n1:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "old";
defparam ram_block1a2.operation_mode = "dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 5;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 31;
defparam ram_block1a2.port_a_logical_ram_depth = 32;
defparam ram_block1a2.port_a_logical_ram_width = 32;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_address_clear = "none";
defparam ram_block1a2.port_b_address_clock = "clock0";
defparam ram_block1a2.port_b_address_width = 5;
defparam ram_block1a2.port_b_data_out_clear = "none";
defparam ram_block1a2.port_b_data_out_clock = "none";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 31;
defparam ram_block1a2.port_b_logical_ram_depth = 32;
defparam ram_block1a2.port_b_logical_ram_width = 32;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock0";
defparam ram_block1a2.ram_block_type = "auto";
defparam ram_block1a2.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a0(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.init_file = "processor_cpu_rf_ram_a.mif";
defparam ram_block1a0.init_file_layout = "port_b";
defparam ram_block1a0.logical_ram_name = "processor_cpu:cpu|processor_cpu_register_bank_a_module:processor_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_44n1:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "old";
defparam ram_block1a0.operation_mode = "dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 5;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 31;
defparam ram_block1a0.port_a_logical_ram_depth = 32;
defparam ram_block1a0.port_a_logical_ram_width = 32;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_address_clear = "none";
defparam ram_block1a0.port_b_address_clock = "clock0";
defparam ram_block1a0.port_b_address_width = 5;
defparam ram_block1a0.port_b_data_out_clear = "none";
defparam ram_block1a0.port_b_data_out_clock = "none";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 31;
defparam ram_block1a0.port_b_logical_ram_depth = 32;
defparam ram_block1a0.port_b_logical_ram_width = 32;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock0";
defparam ram_block1a0.ram_block_type = "auto";
defparam ram_block1a0.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a1(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.init_file = "processor_cpu_rf_ram_a.mif";
defparam ram_block1a1.init_file_layout = "port_b";
defparam ram_block1a1.logical_ram_name = "processor_cpu:cpu|processor_cpu_register_bank_a_module:processor_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_44n1:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "old";
defparam ram_block1a1.operation_mode = "dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 5;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 31;
defparam ram_block1a1.port_a_logical_ram_depth = 32;
defparam ram_block1a1.port_a_logical_ram_width = 32;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_address_clear = "none";
defparam ram_block1a1.port_b_address_clock = "clock0";
defparam ram_block1a1.port_b_address_width = 5;
defparam ram_block1a1.port_b_data_out_clear = "none";
defparam ram_block1a1.port_b_data_out_clock = "none";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 31;
defparam ram_block1a1.port_b_logical_ram_depth = 32;
defparam ram_block1a1.port_b_logical_ram_width = 32;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock0";
defparam ram_block1a1.ram_block_type = "auto";
defparam ram_block1a1.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a31(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[31]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a31_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a31.data_interleave_offset_in_bits = 1;
defparam ram_block1a31.data_interleave_width_in_bits = 1;
defparam ram_block1a31.init_file = "processor_cpu_rf_ram_a.mif";
defparam ram_block1a31.init_file_layout = "port_b";
defparam ram_block1a31.logical_ram_name = "processor_cpu:cpu|processor_cpu_register_bank_a_module:processor_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_44n1:auto_generated|ALTSYNCRAM";
defparam ram_block1a31.mixed_port_feed_through_mode = "old";
defparam ram_block1a31.operation_mode = "dual_port";
defparam ram_block1a31.port_a_address_clear = "none";
defparam ram_block1a31.port_a_address_width = 5;
defparam ram_block1a31.port_a_data_out_clear = "none";
defparam ram_block1a31.port_a_data_out_clock = "none";
defparam ram_block1a31.port_a_data_width = 1;
defparam ram_block1a31.port_a_first_address = 0;
defparam ram_block1a31.port_a_first_bit_number = 31;
defparam ram_block1a31.port_a_last_address = 31;
defparam ram_block1a31.port_a_logical_ram_depth = 32;
defparam ram_block1a31.port_a_logical_ram_width = 32;
defparam ram_block1a31.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a31.port_b_address_clear = "none";
defparam ram_block1a31.port_b_address_clock = "clock0";
defparam ram_block1a31.port_b_address_width = 5;
defparam ram_block1a31.port_b_data_out_clear = "none";
defparam ram_block1a31.port_b_data_out_clock = "none";
defparam ram_block1a31.port_b_data_width = 1;
defparam ram_block1a31.port_b_first_address = 0;
defparam ram_block1a31.port_b_first_bit_number = 31;
defparam ram_block1a31.port_b_last_address = 31;
defparam ram_block1a31.port_b_logical_ram_depth = 32;
defparam ram_block1a31.port_b_logical_ram_width = 32;
defparam ram_block1a31.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a31.port_b_read_enable_clock = "clock0";
defparam ram_block1a31.ram_block_type = "auto";
defparam ram_block1a31.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a17(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[17]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a17_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a17.data_interleave_offset_in_bits = 1;
defparam ram_block1a17.data_interleave_width_in_bits = 1;
defparam ram_block1a17.init_file = "processor_cpu_rf_ram_a.mif";
defparam ram_block1a17.init_file_layout = "port_b";
defparam ram_block1a17.logical_ram_name = "processor_cpu:cpu|processor_cpu_register_bank_a_module:processor_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_44n1:auto_generated|ALTSYNCRAM";
defparam ram_block1a17.mixed_port_feed_through_mode = "old";
defparam ram_block1a17.operation_mode = "dual_port";
defparam ram_block1a17.port_a_address_clear = "none";
defparam ram_block1a17.port_a_address_width = 5;
defparam ram_block1a17.port_a_data_out_clear = "none";
defparam ram_block1a17.port_a_data_out_clock = "none";
defparam ram_block1a17.port_a_data_width = 1;
defparam ram_block1a17.port_a_first_address = 0;
defparam ram_block1a17.port_a_first_bit_number = 17;
defparam ram_block1a17.port_a_last_address = 31;
defparam ram_block1a17.port_a_logical_ram_depth = 32;
defparam ram_block1a17.port_a_logical_ram_width = 32;
defparam ram_block1a17.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a17.port_b_address_clear = "none";
defparam ram_block1a17.port_b_address_clock = "clock0";
defparam ram_block1a17.port_b_address_width = 5;
defparam ram_block1a17.port_b_data_out_clear = "none";
defparam ram_block1a17.port_b_data_out_clock = "none";
defparam ram_block1a17.port_b_data_width = 1;
defparam ram_block1a17.port_b_first_address = 0;
defparam ram_block1a17.port_b_first_bit_number = 17;
defparam ram_block1a17.port_b_last_address = 31;
defparam ram_block1a17.port_b_logical_ram_depth = 32;
defparam ram_block1a17.port_b_logical_ram_width = 32;
defparam ram_block1a17.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a17.port_b_read_enable_clock = "clock0";
defparam ram_block1a17.ram_block_type = "auto";
defparam ram_block1a17.mem_init0 = "00000000";

cyclonev_ram_block ram_block1a30(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[30]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a30_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a30.data_interleave_offset_in_bits = 1;
defparam ram_block1a30.data_interleave_width_in_bits = 1;
defparam ram_block1a30.init_file = "processor_cpu_rf_ram_a.mif";
defparam ram_block1a30.init_file_layout = "port_b";
defparam ram_block1a30.logical_ram_name = "processor_cpu:cpu|processor_cpu_register_bank_a_module:processor_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_44n1:auto_generated|ALTSYNCRAM";
defparam ram_block1a30.mixed_port_feed_through_mode = "old";
defparam ram_block1a30.operation_mode = "dual_port";
defparam ram_block1a30.port_a_address_clear = "none";
defparam ram_block1a30.port_a_address_width = 5;
defparam ram_block1a30.port_a_data_out_clear = "none";
defparam ram_block1a30.port_a_data_out_clock = "none";
defparam ram_block1a30.port_a_data_width = 1;
defparam ram_block1a30.port_a_first_address = 0;
defparam ram_block1a30.port_a_first_bit_number = 30;
defparam ram_block1a30.port_a_last_address = 31;
defparam ram_block1a30.port_a_logical_ram_depth = 32;
defparam ram_block1a30.port_a_logical_ram_width = 32;
defparam ram_block1a30.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a30.port_b_address_clear = "none";
defparam ram_block1a30.port_b_address_clock = "clock0";
defparam ram_block1a30.port_b_address_width = 5;
defparam ram_block1a30.port_b_data_out_clear = "none";
defparam ram_block1a30.port_b_data_out_clock = "none";
defparam ram_block1a30.port_b_data_width = 1;
defparam ram_block1a30.port_b_first_address = 0;
defparam ram_block1a30.port_b_first_bit_number = 30;
defparam ram_block1a30.port_b_last_address = 31;
defparam ram_block1a30.port_b_logical_ram_depth = 32;
defparam ram_block1a30.port_b_logical_ram_width = 32;
defparam ram_block1a30.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a30.port_b_read_enable_clock = "clock0";
defparam ram_block1a30.ram_block_type = "auto";
defparam ram_block1a30.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a18(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[18]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a18_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a18.data_interleave_offset_in_bits = 1;
defparam ram_block1a18.data_interleave_width_in_bits = 1;
defparam ram_block1a18.init_file = "processor_cpu_rf_ram_a.mif";
defparam ram_block1a18.init_file_layout = "port_b";
defparam ram_block1a18.logical_ram_name = "processor_cpu:cpu|processor_cpu_register_bank_a_module:processor_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_44n1:auto_generated|ALTSYNCRAM";
defparam ram_block1a18.mixed_port_feed_through_mode = "old";
defparam ram_block1a18.operation_mode = "dual_port";
defparam ram_block1a18.port_a_address_clear = "none";
defparam ram_block1a18.port_a_address_width = 5;
defparam ram_block1a18.port_a_data_out_clear = "none";
defparam ram_block1a18.port_a_data_out_clock = "none";
defparam ram_block1a18.port_a_data_width = 1;
defparam ram_block1a18.port_a_first_address = 0;
defparam ram_block1a18.port_a_first_bit_number = 18;
defparam ram_block1a18.port_a_last_address = 31;
defparam ram_block1a18.port_a_logical_ram_depth = 32;
defparam ram_block1a18.port_a_logical_ram_width = 32;
defparam ram_block1a18.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a18.port_b_address_clear = "none";
defparam ram_block1a18.port_b_address_clock = "clock0";
defparam ram_block1a18.port_b_address_width = 5;
defparam ram_block1a18.port_b_data_out_clear = "none";
defparam ram_block1a18.port_b_data_out_clock = "none";
defparam ram_block1a18.port_b_data_width = 1;
defparam ram_block1a18.port_b_first_address = 0;
defparam ram_block1a18.port_b_first_bit_number = 18;
defparam ram_block1a18.port_b_last_address = 31;
defparam ram_block1a18.port_b_logical_ram_depth = 32;
defparam ram_block1a18.port_b_logical_ram_width = 32;
defparam ram_block1a18.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a18.port_b_read_enable_clock = "clock0";
defparam ram_block1a18.ram_block_type = "auto";
defparam ram_block1a18.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a29(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[29]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a29_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a29.data_interleave_offset_in_bits = 1;
defparam ram_block1a29.data_interleave_width_in_bits = 1;
defparam ram_block1a29.init_file = "processor_cpu_rf_ram_a.mif";
defparam ram_block1a29.init_file_layout = "port_b";
defparam ram_block1a29.logical_ram_name = "processor_cpu:cpu|processor_cpu_register_bank_a_module:processor_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_44n1:auto_generated|ALTSYNCRAM";
defparam ram_block1a29.mixed_port_feed_through_mode = "old";
defparam ram_block1a29.operation_mode = "dual_port";
defparam ram_block1a29.port_a_address_clear = "none";
defparam ram_block1a29.port_a_address_width = 5;
defparam ram_block1a29.port_a_data_out_clear = "none";
defparam ram_block1a29.port_a_data_out_clock = "none";
defparam ram_block1a29.port_a_data_width = 1;
defparam ram_block1a29.port_a_first_address = 0;
defparam ram_block1a29.port_a_first_bit_number = 29;
defparam ram_block1a29.port_a_last_address = 31;
defparam ram_block1a29.port_a_logical_ram_depth = 32;
defparam ram_block1a29.port_a_logical_ram_width = 32;
defparam ram_block1a29.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a29.port_b_address_clear = "none";
defparam ram_block1a29.port_b_address_clock = "clock0";
defparam ram_block1a29.port_b_address_width = 5;
defparam ram_block1a29.port_b_data_out_clear = "none";
defparam ram_block1a29.port_b_data_out_clock = "none";
defparam ram_block1a29.port_b_data_width = 1;
defparam ram_block1a29.port_b_first_address = 0;
defparam ram_block1a29.port_b_first_bit_number = 29;
defparam ram_block1a29.port_b_last_address = 31;
defparam ram_block1a29.port_b_logical_ram_depth = 32;
defparam ram_block1a29.port_b_logical_ram_width = 32;
defparam ram_block1a29.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a29.port_b_read_enable_clock = "clock0";
defparam ram_block1a29.ram_block_type = "auto";
defparam ram_block1a29.mem_init0 = "00000000";

cyclonev_ram_block ram_block1a19(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[19]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a19_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a19.data_interleave_offset_in_bits = 1;
defparam ram_block1a19.data_interleave_width_in_bits = 1;
defparam ram_block1a19.init_file = "processor_cpu_rf_ram_a.mif";
defparam ram_block1a19.init_file_layout = "port_b";
defparam ram_block1a19.logical_ram_name = "processor_cpu:cpu|processor_cpu_register_bank_a_module:processor_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_44n1:auto_generated|ALTSYNCRAM";
defparam ram_block1a19.mixed_port_feed_through_mode = "old";
defparam ram_block1a19.operation_mode = "dual_port";
defparam ram_block1a19.port_a_address_clear = "none";
defparam ram_block1a19.port_a_address_width = 5;
defparam ram_block1a19.port_a_data_out_clear = "none";
defparam ram_block1a19.port_a_data_out_clock = "none";
defparam ram_block1a19.port_a_data_width = 1;
defparam ram_block1a19.port_a_first_address = 0;
defparam ram_block1a19.port_a_first_bit_number = 19;
defparam ram_block1a19.port_a_last_address = 31;
defparam ram_block1a19.port_a_logical_ram_depth = 32;
defparam ram_block1a19.port_a_logical_ram_width = 32;
defparam ram_block1a19.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a19.port_b_address_clear = "none";
defparam ram_block1a19.port_b_address_clock = "clock0";
defparam ram_block1a19.port_b_address_width = 5;
defparam ram_block1a19.port_b_data_out_clear = "none";
defparam ram_block1a19.port_b_data_out_clock = "none";
defparam ram_block1a19.port_b_data_width = 1;
defparam ram_block1a19.port_b_first_address = 0;
defparam ram_block1a19.port_b_first_bit_number = 19;
defparam ram_block1a19.port_b_last_address = 31;
defparam ram_block1a19.port_b_logical_ram_depth = 32;
defparam ram_block1a19.port_b_logical_ram_width = 32;
defparam ram_block1a19.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a19.port_b_read_enable_clock = "clock0";
defparam ram_block1a19.ram_block_type = "auto";
defparam ram_block1a19.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a28(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[28]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a28_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a28.data_interleave_offset_in_bits = 1;
defparam ram_block1a28.data_interleave_width_in_bits = 1;
defparam ram_block1a28.init_file = "processor_cpu_rf_ram_a.mif";
defparam ram_block1a28.init_file_layout = "port_b";
defparam ram_block1a28.logical_ram_name = "processor_cpu:cpu|processor_cpu_register_bank_a_module:processor_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_44n1:auto_generated|ALTSYNCRAM";
defparam ram_block1a28.mixed_port_feed_through_mode = "old";
defparam ram_block1a28.operation_mode = "dual_port";
defparam ram_block1a28.port_a_address_clear = "none";
defparam ram_block1a28.port_a_address_width = 5;
defparam ram_block1a28.port_a_data_out_clear = "none";
defparam ram_block1a28.port_a_data_out_clock = "none";
defparam ram_block1a28.port_a_data_width = 1;
defparam ram_block1a28.port_a_first_address = 0;
defparam ram_block1a28.port_a_first_bit_number = 28;
defparam ram_block1a28.port_a_last_address = 31;
defparam ram_block1a28.port_a_logical_ram_depth = 32;
defparam ram_block1a28.port_a_logical_ram_width = 32;
defparam ram_block1a28.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a28.port_b_address_clear = "none";
defparam ram_block1a28.port_b_address_clock = "clock0";
defparam ram_block1a28.port_b_address_width = 5;
defparam ram_block1a28.port_b_data_out_clear = "none";
defparam ram_block1a28.port_b_data_out_clock = "none";
defparam ram_block1a28.port_b_data_width = 1;
defparam ram_block1a28.port_b_first_address = 0;
defparam ram_block1a28.port_b_first_bit_number = 28;
defparam ram_block1a28.port_b_last_address = 31;
defparam ram_block1a28.port_b_logical_ram_depth = 32;
defparam ram_block1a28.port_b_logical_ram_width = 32;
defparam ram_block1a28.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a28.port_b_read_enable_clock = "clock0";
defparam ram_block1a28.ram_block_type = "auto";
defparam ram_block1a28.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a24(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[24]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a24_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a24.data_interleave_offset_in_bits = 1;
defparam ram_block1a24.data_interleave_width_in_bits = 1;
defparam ram_block1a24.init_file = "processor_cpu_rf_ram_a.mif";
defparam ram_block1a24.init_file_layout = "port_b";
defparam ram_block1a24.logical_ram_name = "processor_cpu:cpu|processor_cpu_register_bank_a_module:processor_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_44n1:auto_generated|ALTSYNCRAM";
defparam ram_block1a24.mixed_port_feed_through_mode = "old";
defparam ram_block1a24.operation_mode = "dual_port";
defparam ram_block1a24.port_a_address_clear = "none";
defparam ram_block1a24.port_a_address_width = 5;
defparam ram_block1a24.port_a_data_out_clear = "none";
defparam ram_block1a24.port_a_data_out_clock = "none";
defparam ram_block1a24.port_a_data_width = 1;
defparam ram_block1a24.port_a_first_address = 0;
defparam ram_block1a24.port_a_first_bit_number = 24;
defparam ram_block1a24.port_a_last_address = 31;
defparam ram_block1a24.port_a_logical_ram_depth = 32;
defparam ram_block1a24.port_a_logical_ram_width = 32;
defparam ram_block1a24.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a24.port_b_address_clear = "none";
defparam ram_block1a24.port_b_address_clock = "clock0";
defparam ram_block1a24.port_b_address_width = 5;
defparam ram_block1a24.port_b_data_out_clear = "none";
defparam ram_block1a24.port_b_data_out_clock = "none";
defparam ram_block1a24.port_b_data_width = 1;
defparam ram_block1a24.port_b_first_address = 0;
defparam ram_block1a24.port_b_first_bit_number = 24;
defparam ram_block1a24.port_b_last_address = 31;
defparam ram_block1a24.port_b_logical_ram_depth = 32;
defparam ram_block1a24.port_b_logical_ram_width = 32;
defparam ram_block1a24.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a24.port_b_read_enable_clock = "clock0";
defparam ram_block1a24.ram_block_type = "auto";
defparam ram_block1a24.mem_init0 = "00000000";

cyclonev_ram_block ram_block1a21(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[21]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a21_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a21.data_interleave_offset_in_bits = 1;
defparam ram_block1a21.data_interleave_width_in_bits = 1;
defparam ram_block1a21.init_file = "processor_cpu_rf_ram_a.mif";
defparam ram_block1a21.init_file_layout = "port_b";
defparam ram_block1a21.logical_ram_name = "processor_cpu:cpu|processor_cpu_register_bank_a_module:processor_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_44n1:auto_generated|ALTSYNCRAM";
defparam ram_block1a21.mixed_port_feed_through_mode = "old";
defparam ram_block1a21.operation_mode = "dual_port";
defparam ram_block1a21.port_a_address_clear = "none";
defparam ram_block1a21.port_a_address_width = 5;
defparam ram_block1a21.port_a_data_out_clear = "none";
defparam ram_block1a21.port_a_data_out_clock = "none";
defparam ram_block1a21.port_a_data_width = 1;
defparam ram_block1a21.port_a_first_address = 0;
defparam ram_block1a21.port_a_first_bit_number = 21;
defparam ram_block1a21.port_a_last_address = 31;
defparam ram_block1a21.port_a_logical_ram_depth = 32;
defparam ram_block1a21.port_a_logical_ram_width = 32;
defparam ram_block1a21.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a21.port_b_address_clear = "none";
defparam ram_block1a21.port_b_address_clock = "clock0";
defparam ram_block1a21.port_b_address_width = 5;
defparam ram_block1a21.port_b_data_out_clear = "none";
defparam ram_block1a21.port_b_data_out_clock = "none";
defparam ram_block1a21.port_b_data_width = 1;
defparam ram_block1a21.port_b_first_address = 0;
defparam ram_block1a21.port_b_first_bit_number = 21;
defparam ram_block1a21.port_b_last_address = 31;
defparam ram_block1a21.port_b_logical_ram_depth = 32;
defparam ram_block1a21.port_b_logical_ram_width = 32;
defparam ram_block1a21.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a21.port_b_read_enable_clock = "clock0";
defparam ram_block1a21.ram_block_type = "auto";
defparam ram_block1a21.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a20(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[20]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a20_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a20.data_interleave_offset_in_bits = 1;
defparam ram_block1a20.data_interleave_width_in_bits = 1;
defparam ram_block1a20.init_file = "processor_cpu_rf_ram_a.mif";
defparam ram_block1a20.init_file_layout = "port_b";
defparam ram_block1a20.logical_ram_name = "processor_cpu:cpu|processor_cpu_register_bank_a_module:processor_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_44n1:auto_generated|ALTSYNCRAM";
defparam ram_block1a20.mixed_port_feed_through_mode = "old";
defparam ram_block1a20.operation_mode = "dual_port";
defparam ram_block1a20.port_a_address_clear = "none";
defparam ram_block1a20.port_a_address_width = 5;
defparam ram_block1a20.port_a_data_out_clear = "none";
defparam ram_block1a20.port_a_data_out_clock = "none";
defparam ram_block1a20.port_a_data_width = 1;
defparam ram_block1a20.port_a_first_address = 0;
defparam ram_block1a20.port_a_first_bit_number = 20;
defparam ram_block1a20.port_a_last_address = 31;
defparam ram_block1a20.port_a_logical_ram_depth = 32;
defparam ram_block1a20.port_a_logical_ram_width = 32;
defparam ram_block1a20.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a20.port_b_address_clear = "none";
defparam ram_block1a20.port_b_address_clock = "clock0";
defparam ram_block1a20.port_b_address_width = 5;
defparam ram_block1a20.port_b_data_out_clear = "none";
defparam ram_block1a20.port_b_data_out_clock = "none";
defparam ram_block1a20.port_b_data_width = 1;
defparam ram_block1a20.port_b_first_address = 0;
defparam ram_block1a20.port_b_first_bit_number = 20;
defparam ram_block1a20.port_b_last_address = 31;
defparam ram_block1a20.port_b_logical_ram_depth = 32;
defparam ram_block1a20.port_b_logical_ram_width = 32;
defparam ram_block1a20.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a20.port_b_read_enable_clock = "clock0";
defparam ram_block1a20.ram_block_type = "auto";
defparam ram_block1a20.mem_init0 = "00000000";

cyclonev_ram_block ram_block1a22(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[22]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a22_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a22.data_interleave_offset_in_bits = 1;
defparam ram_block1a22.data_interleave_width_in_bits = 1;
defparam ram_block1a22.init_file = "processor_cpu_rf_ram_a.mif";
defparam ram_block1a22.init_file_layout = "port_b";
defparam ram_block1a22.logical_ram_name = "processor_cpu:cpu|processor_cpu_register_bank_a_module:processor_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_44n1:auto_generated|ALTSYNCRAM";
defparam ram_block1a22.mixed_port_feed_through_mode = "old";
defparam ram_block1a22.operation_mode = "dual_port";
defparam ram_block1a22.port_a_address_clear = "none";
defparam ram_block1a22.port_a_address_width = 5;
defparam ram_block1a22.port_a_data_out_clear = "none";
defparam ram_block1a22.port_a_data_out_clock = "none";
defparam ram_block1a22.port_a_data_width = 1;
defparam ram_block1a22.port_a_first_address = 0;
defparam ram_block1a22.port_a_first_bit_number = 22;
defparam ram_block1a22.port_a_last_address = 31;
defparam ram_block1a22.port_a_logical_ram_depth = 32;
defparam ram_block1a22.port_a_logical_ram_width = 32;
defparam ram_block1a22.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a22.port_b_address_clear = "none";
defparam ram_block1a22.port_b_address_clock = "clock0";
defparam ram_block1a22.port_b_address_width = 5;
defparam ram_block1a22.port_b_data_out_clear = "none";
defparam ram_block1a22.port_b_data_out_clock = "none";
defparam ram_block1a22.port_b_data_width = 1;
defparam ram_block1a22.port_b_first_address = 0;
defparam ram_block1a22.port_b_first_bit_number = 22;
defparam ram_block1a22.port_b_last_address = 31;
defparam ram_block1a22.port_b_logical_ram_depth = 32;
defparam ram_block1a22.port_b_logical_ram_width = 32;
defparam ram_block1a22.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a22.port_b_read_enable_clock = "clock0";
defparam ram_block1a22.ram_block_type = "auto";
defparam ram_block1a22.mem_init0 = "00000000";

cyclonev_ram_block ram_block1a23(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[23]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a23_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a23.data_interleave_offset_in_bits = 1;
defparam ram_block1a23.data_interleave_width_in_bits = 1;
defparam ram_block1a23.init_file = "processor_cpu_rf_ram_a.mif";
defparam ram_block1a23.init_file_layout = "port_b";
defparam ram_block1a23.logical_ram_name = "processor_cpu:cpu|processor_cpu_register_bank_a_module:processor_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_44n1:auto_generated|ALTSYNCRAM";
defparam ram_block1a23.mixed_port_feed_through_mode = "old";
defparam ram_block1a23.operation_mode = "dual_port";
defparam ram_block1a23.port_a_address_clear = "none";
defparam ram_block1a23.port_a_address_width = 5;
defparam ram_block1a23.port_a_data_out_clear = "none";
defparam ram_block1a23.port_a_data_out_clock = "none";
defparam ram_block1a23.port_a_data_width = 1;
defparam ram_block1a23.port_a_first_address = 0;
defparam ram_block1a23.port_a_first_bit_number = 23;
defparam ram_block1a23.port_a_last_address = 31;
defparam ram_block1a23.port_a_logical_ram_depth = 32;
defparam ram_block1a23.port_a_logical_ram_width = 32;
defparam ram_block1a23.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a23.port_b_address_clear = "none";
defparam ram_block1a23.port_b_address_clock = "clock0";
defparam ram_block1a23.port_b_address_width = 5;
defparam ram_block1a23.port_b_data_out_clear = "none";
defparam ram_block1a23.port_b_data_out_clock = "none";
defparam ram_block1a23.port_b_data_width = 1;
defparam ram_block1a23.port_b_first_address = 0;
defparam ram_block1a23.port_b_first_bit_number = 23;
defparam ram_block1a23.port_b_last_address = 31;
defparam ram_block1a23.port_b_logical_ram_depth = 32;
defparam ram_block1a23.port_b_logical_ram_width = 32;
defparam ram_block1a23.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a23.port_b_read_enable_clock = "clock0";
defparam ram_block1a23.ram_block_type = "auto";
defparam ram_block1a23.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a27(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[27]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a27_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a27.data_interleave_offset_in_bits = 1;
defparam ram_block1a27.data_interleave_width_in_bits = 1;
defparam ram_block1a27.init_file = "processor_cpu_rf_ram_a.mif";
defparam ram_block1a27.init_file_layout = "port_b";
defparam ram_block1a27.logical_ram_name = "processor_cpu:cpu|processor_cpu_register_bank_a_module:processor_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_44n1:auto_generated|ALTSYNCRAM";
defparam ram_block1a27.mixed_port_feed_through_mode = "old";
defparam ram_block1a27.operation_mode = "dual_port";
defparam ram_block1a27.port_a_address_clear = "none";
defparam ram_block1a27.port_a_address_width = 5;
defparam ram_block1a27.port_a_data_out_clear = "none";
defparam ram_block1a27.port_a_data_out_clock = "none";
defparam ram_block1a27.port_a_data_width = 1;
defparam ram_block1a27.port_a_first_address = 0;
defparam ram_block1a27.port_a_first_bit_number = 27;
defparam ram_block1a27.port_a_last_address = 31;
defparam ram_block1a27.port_a_logical_ram_depth = 32;
defparam ram_block1a27.port_a_logical_ram_width = 32;
defparam ram_block1a27.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a27.port_b_address_clear = "none";
defparam ram_block1a27.port_b_address_clock = "clock0";
defparam ram_block1a27.port_b_address_width = 5;
defparam ram_block1a27.port_b_data_out_clear = "none";
defparam ram_block1a27.port_b_data_out_clock = "none";
defparam ram_block1a27.port_b_data_width = 1;
defparam ram_block1a27.port_b_first_address = 0;
defparam ram_block1a27.port_b_first_bit_number = 27;
defparam ram_block1a27.port_b_last_address = 31;
defparam ram_block1a27.port_b_logical_ram_depth = 32;
defparam ram_block1a27.port_b_logical_ram_width = 32;
defparam ram_block1a27.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a27.port_b_read_enable_clock = "clock0";
defparam ram_block1a27.ram_block_type = "auto";
defparam ram_block1a27.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a26(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[26]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a26_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a26.data_interleave_offset_in_bits = 1;
defparam ram_block1a26.data_interleave_width_in_bits = 1;
defparam ram_block1a26.init_file = "processor_cpu_rf_ram_a.mif";
defparam ram_block1a26.init_file_layout = "port_b";
defparam ram_block1a26.logical_ram_name = "processor_cpu:cpu|processor_cpu_register_bank_a_module:processor_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_44n1:auto_generated|ALTSYNCRAM";
defparam ram_block1a26.mixed_port_feed_through_mode = "old";
defparam ram_block1a26.operation_mode = "dual_port";
defparam ram_block1a26.port_a_address_clear = "none";
defparam ram_block1a26.port_a_address_width = 5;
defparam ram_block1a26.port_a_data_out_clear = "none";
defparam ram_block1a26.port_a_data_out_clock = "none";
defparam ram_block1a26.port_a_data_width = 1;
defparam ram_block1a26.port_a_first_address = 0;
defparam ram_block1a26.port_a_first_bit_number = 26;
defparam ram_block1a26.port_a_last_address = 31;
defparam ram_block1a26.port_a_logical_ram_depth = 32;
defparam ram_block1a26.port_a_logical_ram_width = 32;
defparam ram_block1a26.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a26.port_b_address_clear = "none";
defparam ram_block1a26.port_b_address_clock = "clock0";
defparam ram_block1a26.port_b_address_width = 5;
defparam ram_block1a26.port_b_data_out_clear = "none";
defparam ram_block1a26.port_b_data_out_clock = "none";
defparam ram_block1a26.port_b_data_width = 1;
defparam ram_block1a26.port_b_first_address = 0;
defparam ram_block1a26.port_b_first_bit_number = 26;
defparam ram_block1a26.port_b_last_address = 31;
defparam ram_block1a26.port_b_logical_ram_depth = 32;
defparam ram_block1a26.port_b_logical_ram_width = 32;
defparam ram_block1a26.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a26.port_b_read_enable_clock = "clock0";
defparam ram_block1a26.ram_block_type = "auto";
defparam ram_block1a26.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a25(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[25]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a25_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a25.data_interleave_offset_in_bits = 1;
defparam ram_block1a25.data_interleave_width_in_bits = 1;
defparam ram_block1a25.init_file = "processor_cpu_rf_ram_a.mif";
defparam ram_block1a25.init_file_layout = "port_b";
defparam ram_block1a25.logical_ram_name = "processor_cpu:cpu|processor_cpu_register_bank_a_module:processor_cpu_register_bank_a|altsyncram:the_altsyncram|altsyncram_44n1:auto_generated|ALTSYNCRAM";
defparam ram_block1a25.mixed_port_feed_through_mode = "old";
defparam ram_block1a25.operation_mode = "dual_port";
defparam ram_block1a25.port_a_address_clear = "none";
defparam ram_block1a25.port_a_address_width = 5;
defparam ram_block1a25.port_a_data_out_clear = "none";
defparam ram_block1a25.port_a_data_out_clock = "none";
defparam ram_block1a25.port_a_data_width = 1;
defparam ram_block1a25.port_a_first_address = 0;
defparam ram_block1a25.port_a_first_bit_number = 25;
defparam ram_block1a25.port_a_last_address = 31;
defparam ram_block1a25.port_a_logical_ram_depth = 32;
defparam ram_block1a25.port_a_logical_ram_width = 32;
defparam ram_block1a25.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a25.port_b_address_clear = "none";
defparam ram_block1a25.port_b_address_clock = "clock0";
defparam ram_block1a25.port_b_address_width = 5;
defparam ram_block1a25.port_b_data_out_clear = "none";
defparam ram_block1a25.port_b_data_out_clock = "none";
defparam ram_block1a25.port_b_data_width = 1;
defparam ram_block1a25.port_b_first_address = 0;
defparam ram_block1a25.port_b_first_bit_number = 25;
defparam ram_block1a25.port_b_last_address = 31;
defparam ram_block1a25.port_b_logical_ram_depth = 32;
defparam ram_block1a25.port_b_logical_ram_width = 32;
defparam ram_block1a25.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a25.port_b_read_enable_clock = "clock0";
defparam ram_block1a25.ram_block_type = "auto";
defparam ram_block1a25.mem_init0 = "FFFFFFFF";

endmodule

module processor_processor_cpu_register_bank_b_module (
	q_b_0,
	q_b_5,
	q_b_4,
	q_b_6,
	q_b_16,
	q_b_15,
	q_b_14,
	q_b_13,
	q_b_12,
	q_b_11,
	q_b_10,
	q_b_9,
	q_b_8,
	q_b_7,
	q_b_3,
	q_b_2,
	q_b_1,
	q_b_24,
	q_b_22,
	q_b_23,
	q_b_25,
	q_b_26,
	q_b_31,
	q_b_17,
	q_b_30,
	q_b_241,
	q_b_21,
	q_b_29,
	q_b_20,
	q_b_28,
	q_b_221,
	q_b_18,
	q_b_231,
	q_b_27,
	q_b_261,
	q_b_251,
	q_b_19,
	W_stall,
	M_wr_data_unfiltered_5,
	M_wr_data_unfiltered_15,
	M_wr_data_unfiltered_14,
	M_wr_data_unfiltered_13,
	M_wr_data_unfiltered_12,
	M_wr_data_unfiltered_11,
	M_wr_data_unfiltered_9,
	M_wr_data_unfiltered_7,
	M_wr_data_unfiltered_3,
	M_wr_data_unfiltered_1,
	M_wr_data_unfiltered_0,
	M_dst_regnum_4,
	M_wr_dst_reg,
	M_dst_regnum_0,
	M_dst_regnum_1,
	M_dst_regnum_2,
	M_dst_regnum_3,
	M_wr_data_unfiltered_4,
	M_wr_data_unfiltered_6,
	M_wr_data_unfiltered_16,
	M_wr_data_unfiltered_10,
	M_wr_data_unfiltered_8,
	M_wr_data_unfiltered_2,
	M_wr_data_unfiltered_31,
	M_wr_data_unfiltered_17,
	M_wr_data_unfiltered_30,
	M_wr_data_unfiltered_29,
	M_wr_data_unfiltered_21,
	M_wr_data_unfiltered_19,
	M_wr_data_unfiltered_18,
	M_wr_data_unfiltered_23,
	M_wr_data_unfiltered_27,
	M_wr_data_unfiltered_25,
	M_wr_data_unfiltered_24,
	M_wr_data_unfiltered_20,
	M_wr_data_unfiltered_28,
	M_wr_data_unfiltered_22,
	M_wr_data_unfiltered_26,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_0;
output 	q_b_5;
output 	q_b_4;
output 	q_b_6;
output 	q_b_16;
output 	q_b_15;
output 	q_b_14;
output 	q_b_13;
output 	q_b_12;
output 	q_b_11;
output 	q_b_10;
output 	q_b_9;
output 	q_b_8;
output 	q_b_7;
output 	q_b_3;
output 	q_b_2;
output 	q_b_1;
input 	q_b_24;
input 	q_b_22;
input 	q_b_23;
input 	q_b_25;
input 	q_b_26;
output 	q_b_31;
output 	q_b_17;
output 	q_b_30;
output 	q_b_241;
output 	q_b_21;
output 	q_b_29;
output 	q_b_20;
output 	q_b_28;
output 	q_b_221;
output 	q_b_18;
output 	q_b_231;
output 	q_b_27;
output 	q_b_261;
output 	q_b_251;
output 	q_b_19;
input 	W_stall;
input 	M_wr_data_unfiltered_5;
input 	M_wr_data_unfiltered_15;
input 	M_wr_data_unfiltered_14;
input 	M_wr_data_unfiltered_13;
input 	M_wr_data_unfiltered_12;
input 	M_wr_data_unfiltered_11;
input 	M_wr_data_unfiltered_9;
input 	M_wr_data_unfiltered_7;
input 	M_wr_data_unfiltered_3;
input 	M_wr_data_unfiltered_1;
input 	M_wr_data_unfiltered_0;
input 	M_dst_regnum_4;
input 	M_wr_dst_reg;
input 	M_dst_regnum_0;
input 	M_dst_regnum_1;
input 	M_dst_regnum_2;
input 	M_dst_regnum_3;
input 	M_wr_data_unfiltered_4;
input 	M_wr_data_unfiltered_6;
input 	M_wr_data_unfiltered_16;
input 	M_wr_data_unfiltered_10;
input 	M_wr_data_unfiltered_8;
input 	M_wr_data_unfiltered_2;
input 	M_wr_data_unfiltered_31;
input 	M_wr_data_unfiltered_17;
input 	M_wr_data_unfiltered_30;
input 	M_wr_data_unfiltered_29;
input 	M_wr_data_unfiltered_21;
input 	M_wr_data_unfiltered_19;
input 	M_wr_data_unfiltered_18;
input 	M_wr_data_unfiltered_23;
input 	M_wr_data_unfiltered_27;
input 	M_wr_data_unfiltered_25;
input 	M_wr_data_unfiltered_24;
input 	M_wr_data_unfiltered_20;
input 	M_wr_data_unfiltered_28;
input 	M_wr_data_unfiltered_22;
input 	M_wr_data_unfiltered_26;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



processor_altsyncram_5 the_altsyncram(
	.q_b({q_b_31,q_b_30,q_b_29,q_b_28,q_b_27,q_b_261,q_b_251,q_b_241,q_b_231,q_b_221,q_b_21,q_b_20,q_b_19,q_b_18,q_b_17,q_b_16,q_b_15,q_b_14,q_b_13,q_b_12,q_b_11,q_b_10,q_b_9,q_b_8,q_b_7,q_b_6,q_b_5,q_b_4,q_b_3,q_b_2,q_b_1,q_b_0}),
	.address_b({gnd,gnd,gnd,gnd,q_b_26,q_b_25,q_b_24,q_b_23,q_b_22}),
	.rden_b(W_stall),
	.data_a({M_wr_data_unfiltered_31,M_wr_data_unfiltered_30,M_wr_data_unfiltered_29,M_wr_data_unfiltered_28,M_wr_data_unfiltered_27,M_wr_data_unfiltered_26,M_wr_data_unfiltered_25,M_wr_data_unfiltered_24,M_wr_data_unfiltered_23,M_wr_data_unfiltered_22,M_wr_data_unfiltered_21,
M_wr_data_unfiltered_20,M_wr_data_unfiltered_19,M_wr_data_unfiltered_18,M_wr_data_unfiltered_17,M_wr_data_unfiltered_16,M_wr_data_unfiltered_15,M_wr_data_unfiltered_14,M_wr_data_unfiltered_13,M_wr_data_unfiltered_12,M_wr_data_unfiltered_11,M_wr_data_unfiltered_10,
M_wr_data_unfiltered_9,M_wr_data_unfiltered_8,M_wr_data_unfiltered_7,M_wr_data_unfiltered_6,M_wr_data_unfiltered_5,M_wr_data_unfiltered_4,M_wr_data_unfiltered_3,M_wr_data_unfiltered_2,M_wr_data_unfiltered_1,M_wr_data_unfiltered_0}),
	.address_a({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,M_dst_regnum_4,M_dst_regnum_3,M_dst_regnum_2,M_dst_regnum_1,M_dst_regnum_0}),
	.wren_a(M_wr_dst_reg),
	.clock0(clk_clk));

endmodule

module processor_altsyncram_5 (
	q_b,
	address_b,
	rden_b,
	data_a,
	address_a,
	wren_a,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[31:0] q_b;
input 	[8:0] address_b;
input 	rden_b;
input 	[31:0] data_a;
input 	[12:0] address_a;
input 	wren_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



processor_altsyncram_54n1 auto_generated(
	.q_b({q_b[31],q_b[30],q_b[29],q_b[28],q_b[27],q_b[26],q_b[25],q_b[24],q_b[23],q_b[22],q_b[21],q_b[20],q_b[19],q_b[18],q_b[17],q_b[16],q_b[15],q_b[14],q_b[13],q_b[12],q_b[11],q_b[10],q_b[9],q_b[8],q_b[7],q_b[6],q_b[5],q_b[4],q_b[3],q_b[2],q_b[1],q_b[0]}),
	.address_b({address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.rden_b(rden_b),
	.data_a({data_a[31],data_a[30],data_a[29],data_a[28],data_a[27],data_a[26],data_a[25],data_a[24],data_a[23],data_a[22],data_a[21],data_a[20],data_a[19],data_a[18],data_a[17],data_a[16],data_a[15],data_a[14],data_a[13],data_a[12],data_a[11],data_a[10],data_a[9],data_a[8],data_a[7],data_a[6],data_a[5],data_a[4],data_a[3],data_a[2],data_a[1],data_a[0]}),
	.address_a({address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.wren_a(wren_a),
	.clock0(clock0));

endmodule

module processor_altsyncram_54n1 (
	q_b,
	address_b,
	rden_b,
	data_a,
	address_a,
	wren_a,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[31:0] q_b;
input 	[4:0] address_b;
input 	rden_b;
input 	[31:0] data_a;
input 	[4:0] address_a;
input 	wren_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a0_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a4_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a16_PORTBDATAOUT_bus;
wire [143:0] ram_block1a15_PORTBDATAOUT_bus;
wire [143:0] ram_block1a14_PORTBDATAOUT_bus;
wire [143:0] ram_block1a13_PORTBDATAOUT_bus;
wire [143:0] ram_block1a12_PORTBDATAOUT_bus;
wire [143:0] ram_block1a11_PORTBDATAOUT_bus;
wire [143:0] ram_block1a10_PORTBDATAOUT_bus;
wire [143:0] ram_block1a9_PORTBDATAOUT_bus;
wire [143:0] ram_block1a8_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;
wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a1_PORTBDATAOUT_bus;
wire [143:0] ram_block1a31_PORTBDATAOUT_bus;
wire [143:0] ram_block1a17_PORTBDATAOUT_bus;
wire [143:0] ram_block1a30_PORTBDATAOUT_bus;
wire [143:0] ram_block1a24_PORTBDATAOUT_bus;
wire [143:0] ram_block1a21_PORTBDATAOUT_bus;
wire [143:0] ram_block1a29_PORTBDATAOUT_bus;
wire [143:0] ram_block1a20_PORTBDATAOUT_bus;
wire [143:0] ram_block1a28_PORTBDATAOUT_bus;
wire [143:0] ram_block1a22_PORTBDATAOUT_bus;
wire [143:0] ram_block1a18_PORTBDATAOUT_bus;
wire [143:0] ram_block1a23_PORTBDATAOUT_bus;
wire [143:0] ram_block1a27_PORTBDATAOUT_bus;
wire [143:0] ram_block1a26_PORTBDATAOUT_bus;
wire [143:0] ram_block1a25_PORTBDATAOUT_bus;
wire [143:0] ram_block1a19_PORTBDATAOUT_bus;

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_b[16] = ram_block1a16_PORTBDATAOUT_bus[0];

assign q_b[15] = ram_block1a15_PORTBDATAOUT_bus[0];

assign q_b[14] = ram_block1a14_PORTBDATAOUT_bus[0];

assign q_b[13] = ram_block1a13_PORTBDATAOUT_bus[0];

assign q_b[12] = ram_block1a12_PORTBDATAOUT_bus[0];

assign q_b[11] = ram_block1a11_PORTBDATAOUT_bus[0];

assign q_b[10] = ram_block1a10_PORTBDATAOUT_bus[0];

assign q_b[9] = ram_block1a9_PORTBDATAOUT_bus[0];

assign q_b[8] = ram_block1a8_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_b[3] = ram_block1a3_PORTBDATAOUT_bus[0];

assign q_b[2] = ram_block1a2_PORTBDATAOUT_bus[0];

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

assign q_b[31] = ram_block1a31_PORTBDATAOUT_bus[0];

assign q_b[17] = ram_block1a17_PORTBDATAOUT_bus[0];

assign q_b[30] = ram_block1a30_PORTBDATAOUT_bus[0];

assign q_b[24] = ram_block1a24_PORTBDATAOUT_bus[0];

assign q_b[21] = ram_block1a21_PORTBDATAOUT_bus[0];

assign q_b[29] = ram_block1a29_PORTBDATAOUT_bus[0];

assign q_b[20] = ram_block1a20_PORTBDATAOUT_bus[0];

assign q_b[28] = ram_block1a28_PORTBDATAOUT_bus[0];

assign q_b[22] = ram_block1a22_PORTBDATAOUT_bus[0];

assign q_b[18] = ram_block1a18_PORTBDATAOUT_bus[0];

assign q_b[23] = ram_block1a23_PORTBDATAOUT_bus[0];

assign q_b[27] = ram_block1a27_PORTBDATAOUT_bus[0];

assign q_b[26] = ram_block1a26_PORTBDATAOUT_bus[0];

assign q_b[25] = ram_block1a25_PORTBDATAOUT_bus[0];

assign q_b[19] = ram_block1a19_PORTBDATAOUT_bus[0];

cyclonev_ram_block ram_block1a0(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.init_file = "processor_cpu_rf_ram_b.mif";
defparam ram_block1a0.init_file_layout = "port_b";
defparam ram_block1a0.logical_ram_name = "processor_cpu:cpu|processor_cpu_register_bank_b_module:processor_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_54n1:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "old";
defparam ram_block1a0.operation_mode = "dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 5;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 31;
defparam ram_block1a0.port_a_logical_ram_depth = 32;
defparam ram_block1a0.port_a_logical_ram_width = 32;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_address_clear = "none";
defparam ram_block1a0.port_b_address_clock = "clock0";
defparam ram_block1a0.port_b_address_width = 5;
defparam ram_block1a0.port_b_data_out_clear = "none";
defparam ram_block1a0.port_b_data_out_clock = "none";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 31;
defparam ram_block1a0.port_b_logical_ram_depth = 32;
defparam ram_block1a0.port_b_logical_ram_width = 32;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock0";
defparam ram_block1a0.ram_block_type = "auto";
defparam ram_block1a0.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a5(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.init_file = "processor_cpu_rf_ram_b.mif";
defparam ram_block1a5.init_file_layout = "port_b";
defparam ram_block1a5.logical_ram_name = "processor_cpu:cpu|processor_cpu_register_bank_b_module:processor_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_54n1:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "old";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 5;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 31;
defparam ram_block1a5.port_a_logical_ram_depth = 32;
defparam ram_block1a5.port_a_logical_ram_width = 32;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_address_clear = "none";
defparam ram_block1a5.port_b_address_clock = "clock0";
defparam ram_block1a5.port_b_address_width = 5;
defparam ram_block1a5.port_b_data_out_clear = "none";
defparam ram_block1a5.port_b_data_out_clock = "none";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 31;
defparam ram_block1a5.port_b_logical_ram_depth = 32;
defparam ram_block1a5.port_b_logical_ram_width = 32;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock0";
defparam ram_block1a5.ram_block_type = "auto";
defparam ram_block1a5.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a4(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.init_file = "processor_cpu_rf_ram_b.mif";
defparam ram_block1a4.init_file_layout = "port_b";
defparam ram_block1a4.logical_ram_name = "processor_cpu:cpu|processor_cpu_register_bank_b_module:processor_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_54n1:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "old";
defparam ram_block1a4.operation_mode = "dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 5;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 31;
defparam ram_block1a4.port_a_logical_ram_depth = 32;
defparam ram_block1a4.port_a_logical_ram_width = 32;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_address_clear = "none";
defparam ram_block1a4.port_b_address_clock = "clock0";
defparam ram_block1a4.port_b_address_width = 5;
defparam ram_block1a4.port_b_data_out_clear = "none";
defparam ram_block1a4.port_b_data_out_clock = "none";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 31;
defparam ram_block1a4.port_b_logical_ram_depth = 32;
defparam ram_block1a4.port_b_logical_ram_width = 32;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock0";
defparam ram_block1a4.ram_block_type = "auto";
defparam ram_block1a4.mem_init0 = "00000000";

cyclonev_ram_block ram_block1a6(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.init_file = "processor_cpu_rf_ram_b.mif";
defparam ram_block1a6.init_file_layout = "port_b";
defparam ram_block1a6.logical_ram_name = "processor_cpu:cpu|processor_cpu_register_bank_b_module:processor_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_54n1:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "old";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 5;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 31;
defparam ram_block1a6.port_a_logical_ram_depth = 32;
defparam ram_block1a6.port_a_logical_ram_width = 32;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_address_clear = "none";
defparam ram_block1a6.port_b_address_clock = "clock0";
defparam ram_block1a6.port_b_address_width = 5;
defparam ram_block1a6.port_b_data_out_clear = "none";
defparam ram_block1a6.port_b_data_out_clock = "none";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 31;
defparam ram_block1a6.port_b_logical_ram_depth = 32;
defparam ram_block1a6.port_b_logical_ram_width = 32;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock0";
defparam ram_block1a6.ram_block_type = "auto";
defparam ram_block1a6.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a16(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a16_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a16.data_interleave_offset_in_bits = 1;
defparam ram_block1a16.data_interleave_width_in_bits = 1;
defparam ram_block1a16.init_file = "processor_cpu_rf_ram_b.mif";
defparam ram_block1a16.init_file_layout = "port_b";
defparam ram_block1a16.logical_ram_name = "processor_cpu:cpu|processor_cpu_register_bank_b_module:processor_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_54n1:auto_generated|ALTSYNCRAM";
defparam ram_block1a16.mixed_port_feed_through_mode = "old";
defparam ram_block1a16.operation_mode = "dual_port";
defparam ram_block1a16.port_a_address_clear = "none";
defparam ram_block1a16.port_a_address_width = 5;
defparam ram_block1a16.port_a_data_out_clear = "none";
defparam ram_block1a16.port_a_data_out_clock = "none";
defparam ram_block1a16.port_a_data_width = 1;
defparam ram_block1a16.port_a_first_address = 0;
defparam ram_block1a16.port_a_first_bit_number = 16;
defparam ram_block1a16.port_a_last_address = 31;
defparam ram_block1a16.port_a_logical_ram_depth = 32;
defparam ram_block1a16.port_a_logical_ram_width = 32;
defparam ram_block1a16.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a16.port_b_address_clear = "none";
defparam ram_block1a16.port_b_address_clock = "clock0";
defparam ram_block1a16.port_b_address_width = 5;
defparam ram_block1a16.port_b_data_out_clear = "none";
defparam ram_block1a16.port_b_data_out_clock = "none";
defparam ram_block1a16.port_b_data_width = 1;
defparam ram_block1a16.port_b_first_address = 0;
defparam ram_block1a16.port_b_first_bit_number = 16;
defparam ram_block1a16.port_b_last_address = 31;
defparam ram_block1a16.port_b_logical_ram_depth = 32;
defparam ram_block1a16.port_b_logical_ram_width = 32;
defparam ram_block1a16.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a16.port_b_read_enable_clock = "clock0";
defparam ram_block1a16.ram_block_type = "auto";
defparam ram_block1a16.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a15(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a15_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.init_file = "processor_cpu_rf_ram_b.mif";
defparam ram_block1a15.init_file_layout = "port_b";
defparam ram_block1a15.logical_ram_name = "processor_cpu:cpu|processor_cpu_register_bank_b_module:processor_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_54n1:auto_generated|ALTSYNCRAM";
defparam ram_block1a15.mixed_port_feed_through_mode = "old";
defparam ram_block1a15.operation_mode = "dual_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 5;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 31;
defparam ram_block1a15.port_a_logical_ram_depth = 32;
defparam ram_block1a15.port_a_logical_ram_width = 32;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a15.port_b_address_clear = "none";
defparam ram_block1a15.port_b_address_clock = "clock0";
defparam ram_block1a15.port_b_address_width = 5;
defparam ram_block1a15.port_b_data_out_clear = "none";
defparam ram_block1a15.port_b_data_out_clock = "none";
defparam ram_block1a15.port_b_data_width = 1;
defparam ram_block1a15.port_b_first_address = 0;
defparam ram_block1a15.port_b_first_bit_number = 15;
defparam ram_block1a15.port_b_last_address = 31;
defparam ram_block1a15.port_b_logical_ram_depth = 32;
defparam ram_block1a15.port_b_logical_ram_width = 32;
defparam ram_block1a15.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a15.port_b_read_enable_clock = "clock0";
defparam ram_block1a15.ram_block_type = "auto";
defparam ram_block1a15.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a14(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a14_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.init_file = "processor_cpu_rf_ram_b.mif";
defparam ram_block1a14.init_file_layout = "port_b";
defparam ram_block1a14.logical_ram_name = "processor_cpu:cpu|processor_cpu_register_bank_b_module:processor_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_54n1:auto_generated|ALTSYNCRAM";
defparam ram_block1a14.mixed_port_feed_through_mode = "old";
defparam ram_block1a14.operation_mode = "dual_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 5;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 31;
defparam ram_block1a14.port_a_logical_ram_depth = 32;
defparam ram_block1a14.port_a_logical_ram_width = 32;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a14.port_b_address_clear = "none";
defparam ram_block1a14.port_b_address_clock = "clock0";
defparam ram_block1a14.port_b_address_width = 5;
defparam ram_block1a14.port_b_data_out_clear = "none";
defparam ram_block1a14.port_b_data_out_clock = "none";
defparam ram_block1a14.port_b_data_width = 1;
defparam ram_block1a14.port_b_first_address = 0;
defparam ram_block1a14.port_b_first_bit_number = 14;
defparam ram_block1a14.port_b_last_address = 31;
defparam ram_block1a14.port_b_logical_ram_depth = 32;
defparam ram_block1a14.port_b_logical_ram_width = 32;
defparam ram_block1a14.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a14.port_b_read_enable_clock = "clock0";
defparam ram_block1a14.ram_block_type = "auto";
defparam ram_block1a14.mem_init0 = "00000000";

cyclonev_ram_block ram_block1a13(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a13_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.init_file = "processor_cpu_rf_ram_b.mif";
defparam ram_block1a13.init_file_layout = "port_b";
defparam ram_block1a13.logical_ram_name = "processor_cpu:cpu|processor_cpu_register_bank_b_module:processor_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_54n1:auto_generated|ALTSYNCRAM";
defparam ram_block1a13.mixed_port_feed_through_mode = "old";
defparam ram_block1a13.operation_mode = "dual_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 5;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 31;
defparam ram_block1a13.port_a_logical_ram_depth = 32;
defparam ram_block1a13.port_a_logical_ram_width = 32;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a13.port_b_address_clear = "none";
defparam ram_block1a13.port_b_address_clock = "clock0";
defparam ram_block1a13.port_b_address_width = 5;
defparam ram_block1a13.port_b_data_out_clear = "none";
defparam ram_block1a13.port_b_data_out_clock = "none";
defparam ram_block1a13.port_b_data_width = 1;
defparam ram_block1a13.port_b_first_address = 0;
defparam ram_block1a13.port_b_first_bit_number = 13;
defparam ram_block1a13.port_b_last_address = 31;
defparam ram_block1a13.port_b_logical_ram_depth = 32;
defparam ram_block1a13.port_b_logical_ram_width = 32;
defparam ram_block1a13.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a13.port_b_read_enable_clock = "clock0";
defparam ram_block1a13.ram_block_type = "auto";
defparam ram_block1a13.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a12(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a12_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.init_file = "processor_cpu_rf_ram_b.mif";
defparam ram_block1a12.init_file_layout = "port_b";
defparam ram_block1a12.logical_ram_name = "processor_cpu:cpu|processor_cpu_register_bank_b_module:processor_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_54n1:auto_generated|ALTSYNCRAM";
defparam ram_block1a12.mixed_port_feed_through_mode = "old";
defparam ram_block1a12.operation_mode = "dual_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 5;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 31;
defparam ram_block1a12.port_a_logical_ram_depth = 32;
defparam ram_block1a12.port_a_logical_ram_width = 32;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a12.port_b_address_clear = "none";
defparam ram_block1a12.port_b_address_clock = "clock0";
defparam ram_block1a12.port_b_address_width = 5;
defparam ram_block1a12.port_b_data_out_clear = "none";
defparam ram_block1a12.port_b_data_out_clock = "none";
defparam ram_block1a12.port_b_data_width = 1;
defparam ram_block1a12.port_b_first_address = 0;
defparam ram_block1a12.port_b_first_bit_number = 12;
defparam ram_block1a12.port_b_last_address = 31;
defparam ram_block1a12.port_b_logical_ram_depth = 32;
defparam ram_block1a12.port_b_logical_ram_width = 32;
defparam ram_block1a12.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a12.port_b_read_enable_clock = "clock0";
defparam ram_block1a12.ram_block_type = "auto";
defparam ram_block1a12.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a11(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a11_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.init_file = "processor_cpu_rf_ram_b.mif";
defparam ram_block1a11.init_file_layout = "port_b";
defparam ram_block1a11.logical_ram_name = "processor_cpu:cpu|processor_cpu_register_bank_b_module:processor_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_54n1:auto_generated|ALTSYNCRAM";
defparam ram_block1a11.mixed_port_feed_through_mode = "old";
defparam ram_block1a11.operation_mode = "dual_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 5;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 31;
defparam ram_block1a11.port_a_logical_ram_depth = 32;
defparam ram_block1a11.port_a_logical_ram_width = 32;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a11.port_b_address_clear = "none";
defparam ram_block1a11.port_b_address_clock = "clock0";
defparam ram_block1a11.port_b_address_width = 5;
defparam ram_block1a11.port_b_data_out_clear = "none";
defparam ram_block1a11.port_b_data_out_clock = "none";
defparam ram_block1a11.port_b_data_width = 1;
defparam ram_block1a11.port_b_first_address = 0;
defparam ram_block1a11.port_b_first_bit_number = 11;
defparam ram_block1a11.port_b_last_address = 31;
defparam ram_block1a11.port_b_logical_ram_depth = 32;
defparam ram_block1a11.port_b_logical_ram_width = 32;
defparam ram_block1a11.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a11.port_b_read_enable_clock = "clock0";
defparam ram_block1a11.ram_block_type = "auto";
defparam ram_block1a11.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a10(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a10_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.init_file = "processor_cpu_rf_ram_b.mif";
defparam ram_block1a10.init_file_layout = "port_b";
defparam ram_block1a10.logical_ram_name = "processor_cpu:cpu|processor_cpu_register_bank_b_module:processor_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_54n1:auto_generated|ALTSYNCRAM";
defparam ram_block1a10.mixed_port_feed_through_mode = "old";
defparam ram_block1a10.operation_mode = "dual_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 5;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 31;
defparam ram_block1a10.port_a_logical_ram_depth = 32;
defparam ram_block1a10.port_a_logical_ram_width = 32;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a10.port_b_address_clear = "none";
defparam ram_block1a10.port_b_address_clock = "clock0";
defparam ram_block1a10.port_b_address_width = 5;
defparam ram_block1a10.port_b_data_out_clear = "none";
defparam ram_block1a10.port_b_data_out_clock = "none";
defparam ram_block1a10.port_b_data_width = 1;
defparam ram_block1a10.port_b_first_address = 0;
defparam ram_block1a10.port_b_first_bit_number = 10;
defparam ram_block1a10.port_b_last_address = 31;
defparam ram_block1a10.port_b_logical_ram_depth = 32;
defparam ram_block1a10.port_b_logical_ram_width = 32;
defparam ram_block1a10.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a10.port_b_read_enable_clock = "clock0";
defparam ram_block1a10.ram_block_type = "auto";
defparam ram_block1a10.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a9(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a9_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.init_file = "processor_cpu_rf_ram_b.mif";
defparam ram_block1a9.init_file_layout = "port_b";
defparam ram_block1a9.logical_ram_name = "processor_cpu:cpu|processor_cpu_register_bank_b_module:processor_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_54n1:auto_generated|ALTSYNCRAM";
defparam ram_block1a9.mixed_port_feed_through_mode = "old";
defparam ram_block1a9.operation_mode = "dual_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 5;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 31;
defparam ram_block1a9.port_a_logical_ram_depth = 32;
defparam ram_block1a9.port_a_logical_ram_width = 32;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a9.port_b_address_clear = "none";
defparam ram_block1a9.port_b_address_clock = "clock0";
defparam ram_block1a9.port_b_address_width = 5;
defparam ram_block1a9.port_b_data_out_clear = "none";
defparam ram_block1a9.port_b_data_out_clock = "none";
defparam ram_block1a9.port_b_data_width = 1;
defparam ram_block1a9.port_b_first_address = 0;
defparam ram_block1a9.port_b_first_bit_number = 9;
defparam ram_block1a9.port_b_last_address = 31;
defparam ram_block1a9.port_b_logical_ram_depth = 32;
defparam ram_block1a9.port_b_logical_ram_width = 32;
defparam ram_block1a9.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a9.port_b_read_enable_clock = "clock0";
defparam ram_block1a9.ram_block_type = "auto";
defparam ram_block1a9.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a8(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a8_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.init_file = "processor_cpu_rf_ram_b.mif";
defparam ram_block1a8.init_file_layout = "port_b";
defparam ram_block1a8.logical_ram_name = "processor_cpu:cpu|processor_cpu_register_bank_b_module:processor_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_54n1:auto_generated|ALTSYNCRAM";
defparam ram_block1a8.mixed_port_feed_through_mode = "old";
defparam ram_block1a8.operation_mode = "dual_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 5;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 31;
defparam ram_block1a8.port_a_logical_ram_depth = 32;
defparam ram_block1a8.port_a_logical_ram_width = 32;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a8.port_b_address_clear = "none";
defparam ram_block1a8.port_b_address_clock = "clock0";
defparam ram_block1a8.port_b_address_width = 5;
defparam ram_block1a8.port_b_data_out_clear = "none";
defparam ram_block1a8.port_b_data_out_clock = "none";
defparam ram_block1a8.port_b_data_width = 1;
defparam ram_block1a8.port_b_first_address = 0;
defparam ram_block1a8.port_b_first_bit_number = 8;
defparam ram_block1a8.port_b_last_address = 31;
defparam ram_block1a8.port_b_logical_ram_depth = 32;
defparam ram_block1a8.port_b_logical_ram_width = 32;
defparam ram_block1a8.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a8.port_b_read_enable_clock = "clock0";
defparam ram_block1a8.ram_block_type = "auto";
defparam ram_block1a8.mem_init0 = "00000000";

cyclonev_ram_block ram_block1a7(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.init_file = "processor_cpu_rf_ram_b.mif";
defparam ram_block1a7.init_file_layout = "port_b";
defparam ram_block1a7.logical_ram_name = "processor_cpu:cpu|processor_cpu_register_bank_b_module:processor_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_54n1:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "old";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 5;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 31;
defparam ram_block1a7.port_a_logical_ram_depth = 32;
defparam ram_block1a7.port_a_logical_ram_width = 32;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_address_clear = "none";
defparam ram_block1a7.port_b_address_clock = "clock0";
defparam ram_block1a7.port_b_address_width = 5;
defparam ram_block1a7.port_b_data_out_clear = "none";
defparam ram_block1a7.port_b_data_out_clock = "none";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 31;
defparam ram_block1a7.port_b_logical_ram_depth = 32;
defparam ram_block1a7.port_b_logical_ram_width = 32;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock0";
defparam ram_block1a7.ram_block_type = "auto";
defparam ram_block1a7.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a3(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.init_file = "processor_cpu_rf_ram_b.mif";
defparam ram_block1a3.init_file_layout = "port_b";
defparam ram_block1a3.logical_ram_name = "processor_cpu:cpu|processor_cpu_register_bank_b_module:processor_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_54n1:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "old";
defparam ram_block1a3.operation_mode = "dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 5;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 31;
defparam ram_block1a3.port_a_logical_ram_depth = 32;
defparam ram_block1a3.port_a_logical_ram_width = 32;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_address_clear = "none";
defparam ram_block1a3.port_b_address_clock = "clock0";
defparam ram_block1a3.port_b_address_width = 5;
defparam ram_block1a3.port_b_data_out_clear = "none";
defparam ram_block1a3.port_b_data_out_clock = "none";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 31;
defparam ram_block1a3.port_b_logical_ram_depth = 32;
defparam ram_block1a3.port_b_logical_ram_width = 32;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock0";
defparam ram_block1a3.ram_block_type = "auto";
defparam ram_block1a3.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a2(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.init_file = "processor_cpu_rf_ram_b.mif";
defparam ram_block1a2.init_file_layout = "port_b";
defparam ram_block1a2.logical_ram_name = "processor_cpu:cpu|processor_cpu_register_bank_b_module:processor_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_54n1:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "old";
defparam ram_block1a2.operation_mode = "dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 5;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 31;
defparam ram_block1a2.port_a_logical_ram_depth = 32;
defparam ram_block1a2.port_a_logical_ram_width = 32;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_address_clear = "none";
defparam ram_block1a2.port_b_address_clock = "clock0";
defparam ram_block1a2.port_b_address_width = 5;
defparam ram_block1a2.port_b_data_out_clear = "none";
defparam ram_block1a2.port_b_data_out_clock = "none";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 31;
defparam ram_block1a2.port_b_logical_ram_depth = 32;
defparam ram_block1a2.port_b_logical_ram_width = 32;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock0";
defparam ram_block1a2.ram_block_type = "auto";
defparam ram_block1a2.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a1(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.init_file = "processor_cpu_rf_ram_b.mif";
defparam ram_block1a1.init_file_layout = "port_b";
defparam ram_block1a1.logical_ram_name = "processor_cpu:cpu|processor_cpu_register_bank_b_module:processor_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_54n1:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "old";
defparam ram_block1a1.operation_mode = "dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 5;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 31;
defparam ram_block1a1.port_a_logical_ram_depth = 32;
defparam ram_block1a1.port_a_logical_ram_width = 32;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_address_clear = "none";
defparam ram_block1a1.port_b_address_clock = "clock0";
defparam ram_block1a1.port_b_address_width = 5;
defparam ram_block1a1.port_b_data_out_clear = "none";
defparam ram_block1a1.port_b_data_out_clock = "none";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 31;
defparam ram_block1a1.port_b_logical_ram_depth = 32;
defparam ram_block1a1.port_b_logical_ram_width = 32;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock0";
defparam ram_block1a1.ram_block_type = "auto";
defparam ram_block1a1.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a31(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[31]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a31_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a31.data_interleave_offset_in_bits = 1;
defparam ram_block1a31.data_interleave_width_in_bits = 1;
defparam ram_block1a31.init_file = "processor_cpu_rf_ram_b.mif";
defparam ram_block1a31.init_file_layout = "port_b";
defparam ram_block1a31.logical_ram_name = "processor_cpu:cpu|processor_cpu_register_bank_b_module:processor_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_54n1:auto_generated|ALTSYNCRAM";
defparam ram_block1a31.mixed_port_feed_through_mode = "old";
defparam ram_block1a31.operation_mode = "dual_port";
defparam ram_block1a31.port_a_address_clear = "none";
defparam ram_block1a31.port_a_address_width = 5;
defparam ram_block1a31.port_a_data_out_clear = "none";
defparam ram_block1a31.port_a_data_out_clock = "none";
defparam ram_block1a31.port_a_data_width = 1;
defparam ram_block1a31.port_a_first_address = 0;
defparam ram_block1a31.port_a_first_bit_number = 31;
defparam ram_block1a31.port_a_last_address = 31;
defparam ram_block1a31.port_a_logical_ram_depth = 32;
defparam ram_block1a31.port_a_logical_ram_width = 32;
defparam ram_block1a31.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a31.port_b_address_clear = "none";
defparam ram_block1a31.port_b_address_clock = "clock0";
defparam ram_block1a31.port_b_address_width = 5;
defparam ram_block1a31.port_b_data_out_clear = "none";
defparam ram_block1a31.port_b_data_out_clock = "none";
defparam ram_block1a31.port_b_data_width = 1;
defparam ram_block1a31.port_b_first_address = 0;
defparam ram_block1a31.port_b_first_bit_number = 31;
defparam ram_block1a31.port_b_last_address = 31;
defparam ram_block1a31.port_b_logical_ram_depth = 32;
defparam ram_block1a31.port_b_logical_ram_width = 32;
defparam ram_block1a31.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a31.port_b_read_enable_clock = "clock0";
defparam ram_block1a31.ram_block_type = "auto";
defparam ram_block1a31.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a17(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[17]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a17_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a17.data_interleave_offset_in_bits = 1;
defparam ram_block1a17.data_interleave_width_in_bits = 1;
defparam ram_block1a17.init_file = "processor_cpu_rf_ram_b.mif";
defparam ram_block1a17.init_file_layout = "port_b";
defparam ram_block1a17.logical_ram_name = "processor_cpu:cpu|processor_cpu_register_bank_b_module:processor_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_54n1:auto_generated|ALTSYNCRAM";
defparam ram_block1a17.mixed_port_feed_through_mode = "old";
defparam ram_block1a17.operation_mode = "dual_port";
defparam ram_block1a17.port_a_address_clear = "none";
defparam ram_block1a17.port_a_address_width = 5;
defparam ram_block1a17.port_a_data_out_clear = "none";
defparam ram_block1a17.port_a_data_out_clock = "none";
defparam ram_block1a17.port_a_data_width = 1;
defparam ram_block1a17.port_a_first_address = 0;
defparam ram_block1a17.port_a_first_bit_number = 17;
defparam ram_block1a17.port_a_last_address = 31;
defparam ram_block1a17.port_a_logical_ram_depth = 32;
defparam ram_block1a17.port_a_logical_ram_width = 32;
defparam ram_block1a17.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a17.port_b_address_clear = "none";
defparam ram_block1a17.port_b_address_clock = "clock0";
defparam ram_block1a17.port_b_address_width = 5;
defparam ram_block1a17.port_b_data_out_clear = "none";
defparam ram_block1a17.port_b_data_out_clock = "none";
defparam ram_block1a17.port_b_data_width = 1;
defparam ram_block1a17.port_b_first_address = 0;
defparam ram_block1a17.port_b_first_bit_number = 17;
defparam ram_block1a17.port_b_last_address = 31;
defparam ram_block1a17.port_b_logical_ram_depth = 32;
defparam ram_block1a17.port_b_logical_ram_width = 32;
defparam ram_block1a17.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a17.port_b_read_enable_clock = "clock0";
defparam ram_block1a17.ram_block_type = "auto";
defparam ram_block1a17.mem_init0 = "00000000";

cyclonev_ram_block ram_block1a30(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[30]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a30_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a30.data_interleave_offset_in_bits = 1;
defparam ram_block1a30.data_interleave_width_in_bits = 1;
defparam ram_block1a30.init_file = "processor_cpu_rf_ram_b.mif";
defparam ram_block1a30.init_file_layout = "port_b";
defparam ram_block1a30.logical_ram_name = "processor_cpu:cpu|processor_cpu_register_bank_b_module:processor_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_54n1:auto_generated|ALTSYNCRAM";
defparam ram_block1a30.mixed_port_feed_through_mode = "old";
defparam ram_block1a30.operation_mode = "dual_port";
defparam ram_block1a30.port_a_address_clear = "none";
defparam ram_block1a30.port_a_address_width = 5;
defparam ram_block1a30.port_a_data_out_clear = "none";
defparam ram_block1a30.port_a_data_out_clock = "none";
defparam ram_block1a30.port_a_data_width = 1;
defparam ram_block1a30.port_a_first_address = 0;
defparam ram_block1a30.port_a_first_bit_number = 30;
defparam ram_block1a30.port_a_last_address = 31;
defparam ram_block1a30.port_a_logical_ram_depth = 32;
defparam ram_block1a30.port_a_logical_ram_width = 32;
defparam ram_block1a30.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a30.port_b_address_clear = "none";
defparam ram_block1a30.port_b_address_clock = "clock0";
defparam ram_block1a30.port_b_address_width = 5;
defparam ram_block1a30.port_b_data_out_clear = "none";
defparam ram_block1a30.port_b_data_out_clock = "none";
defparam ram_block1a30.port_b_data_width = 1;
defparam ram_block1a30.port_b_first_address = 0;
defparam ram_block1a30.port_b_first_bit_number = 30;
defparam ram_block1a30.port_b_last_address = 31;
defparam ram_block1a30.port_b_logical_ram_depth = 32;
defparam ram_block1a30.port_b_logical_ram_width = 32;
defparam ram_block1a30.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a30.port_b_read_enable_clock = "clock0";
defparam ram_block1a30.ram_block_type = "auto";
defparam ram_block1a30.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a24(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[24]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a24_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a24.data_interleave_offset_in_bits = 1;
defparam ram_block1a24.data_interleave_width_in_bits = 1;
defparam ram_block1a24.init_file = "processor_cpu_rf_ram_b.mif";
defparam ram_block1a24.init_file_layout = "port_b";
defparam ram_block1a24.logical_ram_name = "processor_cpu:cpu|processor_cpu_register_bank_b_module:processor_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_54n1:auto_generated|ALTSYNCRAM";
defparam ram_block1a24.mixed_port_feed_through_mode = "old";
defparam ram_block1a24.operation_mode = "dual_port";
defparam ram_block1a24.port_a_address_clear = "none";
defparam ram_block1a24.port_a_address_width = 5;
defparam ram_block1a24.port_a_data_out_clear = "none";
defparam ram_block1a24.port_a_data_out_clock = "none";
defparam ram_block1a24.port_a_data_width = 1;
defparam ram_block1a24.port_a_first_address = 0;
defparam ram_block1a24.port_a_first_bit_number = 24;
defparam ram_block1a24.port_a_last_address = 31;
defparam ram_block1a24.port_a_logical_ram_depth = 32;
defparam ram_block1a24.port_a_logical_ram_width = 32;
defparam ram_block1a24.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a24.port_b_address_clear = "none";
defparam ram_block1a24.port_b_address_clock = "clock0";
defparam ram_block1a24.port_b_address_width = 5;
defparam ram_block1a24.port_b_data_out_clear = "none";
defparam ram_block1a24.port_b_data_out_clock = "none";
defparam ram_block1a24.port_b_data_width = 1;
defparam ram_block1a24.port_b_first_address = 0;
defparam ram_block1a24.port_b_first_bit_number = 24;
defparam ram_block1a24.port_b_last_address = 31;
defparam ram_block1a24.port_b_logical_ram_depth = 32;
defparam ram_block1a24.port_b_logical_ram_width = 32;
defparam ram_block1a24.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a24.port_b_read_enable_clock = "clock0";
defparam ram_block1a24.ram_block_type = "auto";
defparam ram_block1a24.mem_init0 = "00000000";

cyclonev_ram_block ram_block1a21(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[21]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a21_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a21.data_interleave_offset_in_bits = 1;
defparam ram_block1a21.data_interleave_width_in_bits = 1;
defparam ram_block1a21.init_file = "processor_cpu_rf_ram_b.mif";
defparam ram_block1a21.init_file_layout = "port_b";
defparam ram_block1a21.logical_ram_name = "processor_cpu:cpu|processor_cpu_register_bank_b_module:processor_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_54n1:auto_generated|ALTSYNCRAM";
defparam ram_block1a21.mixed_port_feed_through_mode = "old";
defparam ram_block1a21.operation_mode = "dual_port";
defparam ram_block1a21.port_a_address_clear = "none";
defparam ram_block1a21.port_a_address_width = 5;
defparam ram_block1a21.port_a_data_out_clear = "none";
defparam ram_block1a21.port_a_data_out_clock = "none";
defparam ram_block1a21.port_a_data_width = 1;
defparam ram_block1a21.port_a_first_address = 0;
defparam ram_block1a21.port_a_first_bit_number = 21;
defparam ram_block1a21.port_a_last_address = 31;
defparam ram_block1a21.port_a_logical_ram_depth = 32;
defparam ram_block1a21.port_a_logical_ram_width = 32;
defparam ram_block1a21.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a21.port_b_address_clear = "none";
defparam ram_block1a21.port_b_address_clock = "clock0";
defparam ram_block1a21.port_b_address_width = 5;
defparam ram_block1a21.port_b_data_out_clear = "none";
defparam ram_block1a21.port_b_data_out_clock = "none";
defparam ram_block1a21.port_b_data_width = 1;
defparam ram_block1a21.port_b_first_address = 0;
defparam ram_block1a21.port_b_first_bit_number = 21;
defparam ram_block1a21.port_b_last_address = 31;
defparam ram_block1a21.port_b_logical_ram_depth = 32;
defparam ram_block1a21.port_b_logical_ram_width = 32;
defparam ram_block1a21.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a21.port_b_read_enable_clock = "clock0";
defparam ram_block1a21.ram_block_type = "auto";
defparam ram_block1a21.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a29(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[29]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a29_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a29.data_interleave_offset_in_bits = 1;
defparam ram_block1a29.data_interleave_width_in_bits = 1;
defparam ram_block1a29.init_file = "processor_cpu_rf_ram_b.mif";
defparam ram_block1a29.init_file_layout = "port_b";
defparam ram_block1a29.logical_ram_name = "processor_cpu:cpu|processor_cpu_register_bank_b_module:processor_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_54n1:auto_generated|ALTSYNCRAM";
defparam ram_block1a29.mixed_port_feed_through_mode = "old";
defparam ram_block1a29.operation_mode = "dual_port";
defparam ram_block1a29.port_a_address_clear = "none";
defparam ram_block1a29.port_a_address_width = 5;
defparam ram_block1a29.port_a_data_out_clear = "none";
defparam ram_block1a29.port_a_data_out_clock = "none";
defparam ram_block1a29.port_a_data_width = 1;
defparam ram_block1a29.port_a_first_address = 0;
defparam ram_block1a29.port_a_first_bit_number = 29;
defparam ram_block1a29.port_a_last_address = 31;
defparam ram_block1a29.port_a_logical_ram_depth = 32;
defparam ram_block1a29.port_a_logical_ram_width = 32;
defparam ram_block1a29.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a29.port_b_address_clear = "none";
defparam ram_block1a29.port_b_address_clock = "clock0";
defparam ram_block1a29.port_b_address_width = 5;
defparam ram_block1a29.port_b_data_out_clear = "none";
defparam ram_block1a29.port_b_data_out_clock = "none";
defparam ram_block1a29.port_b_data_width = 1;
defparam ram_block1a29.port_b_first_address = 0;
defparam ram_block1a29.port_b_first_bit_number = 29;
defparam ram_block1a29.port_b_last_address = 31;
defparam ram_block1a29.port_b_logical_ram_depth = 32;
defparam ram_block1a29.port_b_logical_ram_width = 32;
defparam ram_block1a29.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a29.port_b_read_enable_clock = "clock0";
defparam ram_block1a29.ram_block_type = "auto";
defparam ram_block1a29.mem_init0 = "00000000";

cyclonev_ram_block ram_block1a20(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[20]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a20_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a20.data_interleave_offset_in_bits = 1;
defparam ram_block1a20.data_interleave_width_in_bits = 1;
defparam ram_block1a20.init_file = "processor_cpu_rf_ram_b.mif";
defparam ram_block1a20.init_file_layout = "port_b";
defparam ram_block1a20.logical_ram_name = "processor_cpu:cpu|processor_cpu_register_bank_b_module:processor_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_54n1:auto_generated|ALTSYNCRAM";
defparam ram_block1a20.mixed_port_feed_through_mode = "old";
defparam ram_block1a20.operation_mode = "dual_port";
defparam ram_block1a20.port_a_address_clear = "none";
defparam ram_block1a20.port_a_address_width = 5;
defparam ram_block1a20.port_a_data_out_clear = "none";
defparam ram_block1a20.port_a_data_out_clock = "none";
defparam ram_block1a20.port_a_data_width = 1;
defparam ram_block1a20.port_a_first_address = 0;
defparam ram_block1a20.port_a_first_bit_number = 20;
defparam ram_block1a20.port_a_last_address = 31;
defparam ram_block1a20.port_a_logical_ram_depth = 32;
defparam ram_block1a20.port_a_logical_ram_width = 32;
defparam ram_block1a20.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a20.port_b_address_clear = "none";
defparam ram_block1a20.port_b_address_clock = "clock0";
defparam ram_block1a20.port_b_address_width = 5;
defparam ram_block1a20.port_b_data_out_clear = "none";
defparam ram_block1a20.port_b_data_out_clock = "none";
defparam ram_block1a20.port_b_data_width = 1;
defparam ram_block1a20.port_b_first_address = 0;
defparam ram_block1a20.port_b_first_bit_number = 20;
defparam ram_block1a20.port_b_last_address = 31;
defparam ram_block1a20.port_b_logical_ram_depth = 32;
defparam ram_block1a20.port_b_logical_ram_width = 32;
defparam ram_block1a20.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a20.port_b_read_enable_clock = "clock0";
defparam ram_block1a20.ram_block_type = "auto";
defparam ram_block1a20.mem_init0 = "00000000";

cyclonev_ram_block ram_block1a28(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[28]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a28_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a28.data_interleave_offset_in_bits = 1;
defparam ram_block1a28.data_interleave_width_in_bits = 1;
defparam ram_block1a28.init_file = "processor_cpu_rf_ram_b.mif";
defparam ram_block1a28.init_file_layout = "port_b";
defparam ram_block1a28.logical_ram_name = "processor_cpu:cpu|processor_cpu_register_bank_b_module:processor_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_54n1:auto_generated|ALTSYNCRAM";
defparam ram_block1a28.mixed_port_feed_through_mode = "old";
defparam ram_block1a28.operation_mode = "dual_port";
defparam ram_block1a28.port_a_address_clear = "none";
defparam ram_block1a28.port_a_address_width = 5;
defparam ram_block1a28.port_a_data_out_clear = "none";
defparam ram_block1a28.port_a_data_out_clock = "none";
defparam ram_block1a28.port_a_data_width = 1;
defparam ram_block1a28.port_a_first_address = 0;
defparam ram_block1a28.port_a_first_bit_number = 28;
defparam ram_block1a28.port_a_last_address = 31;
defparam ram_block1a28.port_a_logical_ram_depth = 32;
defparam ram_block1a28.port_a_logical_ram_width = 32;
defparam ram_block1a28.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a28.port_b_address_clear = "none";
defparam ram_block1a28.port_b_address_clock = "clock0";
defparam ram_block1a28.port_b_address_width = 5;
defparam ram_block1a28.port_b_data_out_clear = "none";
defparam ram_block1a28.port_b_data_out_clock = "none";
defparam ram_block1a28.port_b_data_width = 1;
defparam ram_block1a28.port_b_first_address = 0;
defparam ram_block1a28.port_b_first_bit_number = 28;
defparam ram_block1a28.port_b_last_address = 31;
defparam ram_block1a28.port_b_logical_ram_depth = 32;
defparam ram_block1a28.port_b_logical_ram_width = 32;
defparam ram_block1a28.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a28.port_b_read_enable_clock = "clock0";
defparam ram_block1a28.ram_block_type = "auto";
defparam ram_block1a28.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a22(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[22]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a22_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a22.data_interleave_offset_in_bits = 1;
defparam ram_block1a22.data_interleave_width_in_bits = 1;
defparam ram_block1a22.init_file = "processor_cpu_rf_ram_b.mif";
defparam ram_block1a22.init_file_layout = "port_b";
defparam ram_block1a22.logical_ram_name = "processor_cpu:cpu|processor_cpu_register_bank_b_module:processor_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_54n1:auto_generated|ALTSYNCRAM";
defparam ram_block1a22.mixed_port_feed_through_mode = "old";
defparam ram_block1a22.operation_mode = "dual_port";
defparam ram_block1a22.port_a_address_clear = "none";
defparam ram_block1a22.port_a_address_width = 5;
defparam ram_block1a22.port_a_data_out_clear = "none";
defparam ram_block1a22.port_a_data_out_clock = "none";
defparam ram_block1a22.port_a_data_width = 1;
defparam ram_block1a22.port_a_first_address = 0;
defparam ram_block1a22.port_a_first_bit_number = 22;
defparam ram_block1a22.port_a_last_address = 31;
defparam ram_block1a22.port_a_logical_ram_depth = 32;
defparam ram_block1a22.port_a_logical_ram_width = 32;
defparam ram_block1a22.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a22.port_b_address_clear = "none";
defparam ram_block1a22.port_b_address_clock = "clock0";
defparam ram_block1a22.port_b_address_width = 5;
defparam ram_block1a22.port_b_data_out_clear = "none";
defparam ram_block1a22.port_b_data_out_clock = "none";
defparam ram_block1a22.port_b_data_width = 1;
defparam ram_block1a22.port_b_first_address = 0;
defparam ram_block1a22.port_b_first_bit_number = 22;
defparam ram_block1a22.port_b_last_address = 31;
defparam ram_block1a22.port_b_logical_ram_depth = 32;
defparam ram_block1a22.port_b_logical_ram_width = 32;
defparam ram_block1a22.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a22.port_b_read_enable_clock = "clock0";
defparam ram_block1a22.ram_block_type = "auto";
defparam ram_block1a22.mem_init0 = "00000000";

cyclonev_ram_block ram_block1a18(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[18]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a18_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a18.data_interleave_offset_in_bits = 1;
defparam ram_block1a18.data_interleave_width_in_bits = 1;
defparam ram_block1a18.init_file = "processor_cpu_rf_ram_b.mif";
defparam ram_block1a18.init_file_layout = "port_b";
defparam ram_block1a18.logical_ram_name = "processor_cpu:cpu|processor_cpu_register_bank_b_module:processor_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_54n1:auto_generated|ALTSYNCRAM";
defparam ram_block1a18.mixed_port_feed_through_mode = "old";
defparam ram_block1a18.operation_mode = "dual_port";
defparam ram_block1a18.port_a_address_clear = "none";
defparam ram_block1a18.port_a_address_width = 5;
defparam ram_block1a18.port_a_data_out_clear = "none";
defparam ram_block1a18.port_a_data_out_clock = "none";
defparam ram_block1a18.port_a_data_width = 1;
defparam ram_block1a18.port_a_first_address = 0;
defparam ram_block1a18.port_a_first_bit_number = 18;
defparam ram_block1a18.port_a_last_address = 31;
defparam ram_block1a18.port_a_logical_ram_depth = 32;
defparam ram_block1a18.port_a_logical_ram_width = 32;
defparam ram_block1a18.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a18.port_b_address_clear = "none";
defparam ram_block1a18.port_b_address_clock = "clock0";
defparam ram_block1a18.port_b_address_width = 5;
defparam ram_block1a18.port_b_data_out_clear = "none";
defparam ram_block1a18.port_b_data_out_clock = "none";
defparam ram_block1a18.port_b_data_width = 1;
defparam ram_block1a18.port_b_first_address = 0;
defparam ram_block1a18.port_b_first_bit_number = 18;
defparam ram_block1a18.port_b_last_address = 31;
defparam ram_block1a18.port_b_logical_ram_depth = 32;
defparam ram_block1a18.port_b_logical_ram_width = 32;
defparam ram_block1a18.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a18.port_b_read_enable_clock = "clock0";
defparam ram_block1a18.ram_block_type = "auto";
defparam ram_block1a18.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a23(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[23]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a23_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a23.data_interleave_offset_in_bits = 1;
defparam ram_block1a23.data_interleave_width_in_bits = 1;
defparam ram_block1a23.init_file = "processor_cpu_rf_ram_b.mif";
defparam ram_block1a23.init_file_layout = "port_b";
defparam ram_block1a23.logical_ram_name = "processor_cpu:cpu|processor_cpu_register_bank_b_module:processor_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_54n1:auto_generated|ALTSYNCRAM";
defparam ram_block1a23.mixed_port_feed_through_mode = "old";
defparam ram_block1a23.operation_mode = "dual_port";
defparam ram_block1a23.port_a_address_clear = "none";
defparam ram_block1a23.port_a_address_width = 5;
defparam ram_block1a23.port_a_data_out_clear = "none";
defparam ram_block1a23.port_a_data_out_clock = "none";
defparam ram_block1a23.port_a_data_width = 1;
defparam ram_block1a23.port_a_first_address = 0;
defparam ram_block1a23.port_a_first_bit_number = 23;
defparam ram_block1a23.port_a_last_address = 31;
defparam ram_block1a23.port_a_logical_ram_depth = 32;
defparam ram_block1a23.port_a_logical_ram_width = 32;
defparam ram_block1a23.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a23.port_b_address_clear = "none";
defparam ram_block1a23.port_b_address_clock = "clock0";
defparam ram_block1a23.port_b_address_width = 5;
defparam ram_block1a23.port_b_data_out_clear = "none";
defparam ram_block1a23.port_b_data_out_clock = "none";
defparam ram_block1a23.port_b_data_width = 1;
defparam ram_block1a23.port_b_first_address = 0;
defparam ram_block1a23.port_b_first_bit_number = 23;
defparam ram_block1a23.port_b_last_address = 31;
defparam ram_block1a23.port_b_logical_ram_depth = 32;
defparam ram_block1a23.port_b_logical_ram_width = 32;
defparam ram_block1a23.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a23.port_b_read_enable_clock = "clock0";
defparam ram_block1a23.ram_block_type = "auto";
defparam ram_block1a23.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a27(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[27]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a27_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a27.data_interleave_offset_in_bits = 1;
defparam ram_block1a27.data_interleave_width_in_bits = 1;
defparam ram_block1a27.init_file = "processor_cpu_rf_ram_b.mif";
defparam ram_block1a27.init_file_layout = "port_b";
defparam ram_block1a27.logical_ram_name = "processor_cpu:cpu|processor_cpu_register_bank_b_module:processor_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_54n1:auto_generated|ALTSYNCRAM";
defparam ram_block1a27.mixed_port_feed_through_mode = "old";
defparam ram_block1a27.operation_mode = "dual_port";
defparam ram_block1a27.port_a_address_clear = "none";
defparam ram_block1a27.port_a_address_width = 5;
defparam ram_block1a27.port_a_data_out_clear = "none";
defparam ram_block1a27.port_a_data_out_clock = "none";
defparam ram_block1a27.port_a_data_width = 1;
defparam ram_block1a27.port_a_first_address = 0;
defparam ram_block1a27.port_a_first_bit_number = 27;
defparam ram_block1a27.port_a_last_address = 31;
defparam ram_block1a27.port_a_logical_ram_depth = 32;
defparam ram_block1a27.port_a_logical_ram_width = 32;
defparam ram_block1a27.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a27.port_b_address_clear = "none";
defparam ram_block1a27.port_b_address_clock = "clock0";
defparam ram_block1a27.port_b_address_width = 5;
defparam ram_block1a27.port_b_data_out_clear = "none";
defparam ram_block1a27.port_b_data_out_clock = "none";
defparam ram_block1a27.port_b_data_width = 1;
defparam ram_block1a27.port_b_first_address = 0;
defparam ram_block1a27.port_b_first_bit_number = 27;
defparam ram_block1a27.port_b_last_address = 31;
defparam ram_block1a27.port_b_logical_ram_depth = 32;
defparam ram_block1a27.port_b_logical_ram_width = 32;
defparam ram_block1a27.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a27.port_b_read_enable_clock = "clock0";
defparam ram_block1a27.ram_block_type = "auto";
defparam ram_block1a27.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a26(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[26]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a26_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a26.data_interleave_offset_in_bits = 1;
defparam ram_block1a26.data_interleave_width_in_bits = 1;
defparam ram_block1a26.init_file = "processor_cpu_rf_ram_b.mif";
defparam ram_block1a26.init_file_layout = "port_b";
defparam ram_block1a26.logical_ram_name = "processor_cpu:cpu|processor_cpu_register_bank_b_module:processor_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_54n1:auto_generated|ALTSYNCRAM";
defparam ram_block1a26.mixed_port_feed_through_mode = "old";
defparam ram_block1a26.operation_mode = "dual_port";
defparam ram_block1a26.port_a_address_clear = "none";
defparam ram_block1a26.port_a_address_width = 5;
defparam ram_block1a26.port_a_data_out_clear = "none";
defparam ram_block1a26.port_a_data_out_clock = "none";
defparam ram_block1a26.port_a_data_width = 1;
defparam ram_block1a26.port_a_first_address = 0;
defparam ram_block1a26.port_a_first_bit_number = 26;
defparam ram_block1a26.port_a_last_address = 31;
defparam ram_block1a26.port_a_logical_ram_depth = 32;
defparam ram_block1a26.port_a_logical_ram_width = 32;
defparam ram_block1a26.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a26.port_b_address_clear = "none";
defparam ram_block1a26.port_b_address_clock = "clock0";
defparam ram_block1a26.port_b_address_width = 5;
defparam ram_block1a26.port_b_data_out_clear = "none";
defparam ram_block1a26.port_b_data_out_clock = "none";
defparam ram_block1a26.port_b_data_width = 1;
defparam ram_block1a26.port_b_first_address = 0;
defparam ram_block1a26.port_b_first_bit_number = 26;
defparam ram_block1a26.port_b_last_address = 31;
defparam ram_block1a26.port_b_logical_ram_depth = 32;
defparam ram_block1a26.port_b_logical_ram_width = 32;
defparam ram_block1a26.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a26.port_b_read_enable_clock = "clock0";
defparam ram_block1a26.ram_block_type = "auto";
defparam ram_block1a26.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a25(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[25]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a25_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a25.data_interleave_offset_in_bits = 1;
defparam ram_block1a25.data_interleave_width_in_bits = 1;
defparam ram_block1a25.init_file = "processor_cpu_rf_ram_b.mif";
defparam ram_block1a25.init_file_layout = "port_b";
defparam ram_block1a25.logical_ram_name = "processor_cpu:cpu|processor_cpu_register_bank_b_module:processor_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_54n1:auto_generated|ALTSYNCRAM";
defparam ram_block1a25.mixed_port_feed_through_mode = "old";
defparam ram_block1a25.operation_mode = "dual_port";
defparam ram_block1a25.port_a_address_clear = "none";
defparam ram_block1a25.port_a_address_width = 5;
defparam ram_block1a25.port_a_data_out_clear = "none";
defparam ram_block1a25.port_a_data_out_clock = "none";
defparam ram_block1a25.port_a_data_width = 1;
defparam ram_block1a25.port_a_first_address = 0;
defparam ram_block1a25.port_a_first_bit_number = 25;
defparam ram_block1a25.port_a_last_address = 31;
defparam ram_block1a25.port_a_logical_ram_depth = 32;
defparam ram_block1a25.port_a_logical_ram_width = 32;
defparam ram_block1a25.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a25.port_b_address_clear = "none";
defparam ram_block1a25.port_b_address_clock = "clock0";
defparam ram_block1a25.port_b_address_width = 5;
defparam ram_block1a25.port_b_data_out_clear = "none";
defparam ram_block1a25.port_b_data_out_clock = "none";
defparam ram_block1a25.port_b_data_width = 1;
defparam ram_block1a25.port_b_first_address = 0;
defparam ram_block1a25.port_b_first_bit_number = 25;
defparam ram_block1a25.port_b_last_address = 31;
defparam ram_block1a25.port_b_logical_ram_depth = 32;
defparam ram_block1a25.port_b_logical_ram_width = 32;
defparam ram_block1a25.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a25.port_b_read_enable_clock = "clock0";
defparam ram_block1a25.ram_block_type = "auto";
defparam ram_block1a25.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a19(
	.portawe(!wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[19]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a19_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a19.data_interleave_offset_in_bits = 1;
defparam ram_block1a19.data_interleave_width_in_bits = 1;
defparam ram_block1a19.init_file = "processor_cpu_rf_ram_b.mif";
defparam ram_block1a19.init_file_layout = "port_b";
defparam ram_block1a19.logical_ram_name = "processor_cpu:cpu|processor_cpu_register_bank_b_module:processor_cpu_register_bank_b|altsyncram:the_altsyncram|altsyncram_54n1:auto_generated|ALTSYNCRAM";
defparam ram_block1a19.mixed_port_feed_through_mode = "old";
defparam ram_block1a19.operation_mode = "dual_port";
defparam ram_block1a19.port_a_address_clear = "none";
defparam ram_block1a19.port_a_address_width = 5;
defparam ram_block1a19.port_a_data_out_clear = "none";
defparam ram_block1a19.port_a_data_out_clock = "none";
defparam ram_block1a19.port_a_data_width = 1;
defparam ram_block1a19.port_a_first_address = 0;
defparam ram_block1a19.port_a_first_bit_number = 19;
defparam ram_block1a19.port_a_last_address = 31;
defparam ram_block1a19.port_a_logical_ram_depth = 32;
defparam ram_block1a19.port_a_logical_ram_width = 32;
defparam ram_block1a19.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a19.port_b_address_clear = "none";
defparam ram_block1a19.port_b_address_clock = "clock0";
defparam ram_block1a19.port_b_address_width = 5;
defparam ram_block1a19.port_b_data_out_clear = "none";
defparam ram_block1a19.port_b_data_out_clock = "none";
defparam ram_block1a19.port_b_data_width = 1;
defparam ram_block1a19.port_b_first_address = 0;
defparam ram_block1a19.port_b_first_bit_number = 19;
defparam ram_block1a19.port_b_last_address = 31;
defparam ram_block1a19.port_b_logical_ram_depth = 32;
defparam ram_block1a19.port_b_logical_ram_width = 32;
defparam ram_block1a19.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a19.port_b_read_enable_clock = "clock0";
defparam ram_block1a19.ram_block_type = "auto";
defparam ram_block1a19.mem_init0 = "FFFFFFFF";

endmodule

module processor_processor_jtag_uart (
	q_b_0,
	Add1,
	q_b_5,
	Add11,
	q_b_4,
	Add12,
	q_b_6,
	Add13,
	q_b_7,
	M_st_data_10,
	q_b_3,
	Add14,
	q_b_2,
	Add15,
	q_b_1,
	Add16,
	tdo,
	M_st_data_0,
	r_sync_rst,
	clr_break_line,
	d_write,
	Equal1,
	Equal2,
	M_alu_result_2,
	M_st_data_1,
	M_st_data_2,
	M_st_data_3,
	M_st_data_4,
	M_st_data_5,
	M_st_data_6,
	M_st_data_7,
	d_read,
	read_accepted,
	av_waitrequest1,
	Equal6,
	uav_read,
	read_latency_shift_reg,
	ien_AE1,
	av_readdata_9,
	ien_AF1,
	av_readdata_8,
	b_full,
	read_01,
	counter_reg_bit_0,
	counter_reg_bit_5,
	b_full1,
	counter_reg_bit_4,
	b_non_empty,
	woverflow1,
	rvalid1,
	ac1,
	counter_reg_bit_3,
	counter_reg_bit_2,
	counter_reg_bit_1,
	altera_internal_jtag,
	altera_internal_jtag1,
	state_4,
	splitter_nodes_receive_0_3,
	virtual_ir_scan_reg,
	clr_reg,
	state_3,
	state_8,
	irf_reg_0_1,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_0;
output 	Add1;
output 	q_b_5;
output 	Add11;
output 	q_b_4;
output 	Add12;
output 	q_b_6;
output 	Add13;
output 	q_b_7;
input 	M_st_data_10;
output 	q_b_3;
output 	Add14;
output 	q_b_2;
output 	Add15;
output 	q_b_1;
output 	Add16;
output 	tdo;
input 	M_st_data_0;
input 	r_sync_rst;
input 	clr_break_line;
input 	d_write;
input 	Equal1;
input 	Equal2;
input 	M_alu_result_2;
input 	M_st_data_1;
input 	M_st_data_2;
input 	M_st_data_3;
input 	M_st_data_4;
input 	M_st_data_5;
input 	M_st_data_6;
input 	M_st_data_7;
input 	d_read;
input 	read_accepted;
output 	av_waitrequest1;
input 	Equal6;
input 	uav_read;
input 	read_latency_shift_reg;
output 	ien_AE1;
output 	av_readdata_9;
output 	ien_AF1;
output 	av_readdata_8;
output 	b_full;
output 	read_01;
output 	counter_reg_bit_0;
output 	counter_reg_bit_5;
output 	b_full1;
output 	counter_reg_bit_4;
output 	b_non_empty;
output 	woverflow1;
output 	rvalid1;
output 	ac1;
output 	counter_reg_bit_3;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
input 	altera_internal_jtag;
input 	altera_internal_jtag1;
input 	state_4;
input 	splitter_nodes_receive_0_3;
input 	virtual_ir_scan_reg;
input 	clr_reg;
input 	state_3;
input 	state_8;
input 	irf_reg_0_1;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \the_processor_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[7] ;
wire \the_processor_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[0] ;
wire \the_processor_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[1] ;
wire \the_processor_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[2] ;
wire \the_processor_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[3] ;
wire \the_processor_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[6] ;
wire \the_processor_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[5] ;
wire \the_processor_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[4] ;
wire \t_dav~q ;
wire \r_val~q ;
wire \the_processor_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[5]~q ;
wire \the_processor_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[4]~q ;
wire \the_processor_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[0]~q ;
wire \the_processor_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[3]~q ;
wire \the_processor_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[2]~q ;
wire \the_processor_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[1]~q ;
wire \processor_jtag_uart_alt_jtag_atlantic|t_pause~q ;
wire \fifo_wr~q ;
wire \processor_jtag_uart_alt_jtag_atlantic|rvalid0~1_combout ;
wire \the_processor_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|b_non_empty~q ;
wire \r_val~0_combout ;
wire \fifo_rd~2_combout ;
wire \processor_jtag_uart_alt_jtag_atlantic|t_ena~q ;
wire \wr_rfifo~combout ;
wire \processor_jtag_uart_alt_jtag_atlantic|wdata[0]~q ;
wire \processor_jtag_uart_alt_jtag_atlantic|wdata[5]~q ;
wire \processor_jtag_uart_alt_jtag_atlantic|wdata[4]~q ;
wire \processor_jtag_uart_alt_jtag_atlantic|wdata[6]~q ;
wire \processor_jtag_uart_alt_jtag_atlantic|wdata[7]~q ;
wire \processor_jtag_uart_alt_jtag_atlantic|wdata[3]~q ;
wire \processor_jtag_uart_alt_jtag_atlantic|wdata[2]~q ;
wire \processor_jtag_uart_alt_jtag_atlantic|wdata[1]~q ;
wire \fifo_wr~0_combout ;
wire \Add1~2 ;
wire \Add1~6 ;
wire \Add1~10 ;
wire \Add1~18 ;
wire \Add1~22 ;
wire \Add1~26 ;
wire \av_waitrequest~0_combout ;
wire \av_waitrequest~1_combout ;
wire \ien_AE~0_combout ;
wire \LessThan0~0_combout ;
wire \LessThan0~1_combout ;
wire \fifo_AE~q ;
wire \pause_irq~0_combout ;
wire \pause_irq~q ;
wire \Add0~22 ;
wire \Add0~26 ;
wire \Add0~18 ;
wire \Add0~1_sumout ;
wire \Add0~2 ;
wire \Add0~5_sumout ;
wire \Add0~6 ;
wire \Add0~9_sumout ;
wire \Add0~10 ;
wire \Add0~13_sumout ;
wire \Add0~17_sumout ;
wire \Add0~21_sumout ;
wire \Add0~25_sumout ;
wire \LessThan1~0_combout ;
wire \LessThan1~1_combout ;
wire \fifo_AF~q ;
wire \fifo_rd~0_combout ;
wire \fifo_rd~1_combout ;
wire \woverflow~0_combout ;
wire \rvalid~0_combout ;
wire \ac~0_combout ;


processor_processor_jtag_uart_scfifo_w the_processor_jtag_uart_scfifo_w(
	.q_b_7(\the_processor_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[7] ),
	.q_b_0(\the_processor_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[0] ),
	.q_b_1(\the_processor_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[1] ),
	.q_b_2(\the_processor_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[2] ),
	.q_b_3(\the_processor_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[3] ),
	.q_b_6(\the_processor_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[6] ),
	.q_b_5(\the_processor_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[5] ),
	.q_b_4(\the_processor_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[4] ),
	.M_st_data_0(M_st_data_0),
	.r_sync_rst(r_sync_rst),
	.M_st_data_1(M_st_data_1),
	.M_st_data_2(M_st_data_2),
	.M_st_data_3(M_st_data_3),
	.M_st_data_4(M_st_data_4),
	.M_st_data_5(M_st_data_5),
	.M_st_data_6(M_st_data_6),
	.M_st_data_7(M_st_data_7),
	.b_full(b_full1),
	.counter_reg_bit_5(\the_processor_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[5]~q ),
	.counter_reg_bit_4(\the_processor_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[4]~q ),
	.counter_reg_bit_0(\the_processor_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[0]~q ),
	.counter_reg_bit_3(\the_processor_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[3]~q ),
	.counter_reg_bit_2(\the_processor_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[2]~q ),
	.counter_reg_bit_1(\the_processor_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[1]~q ),
	.fifo_wr(\fifo_wr~q ),
	.b_non_empty(\the_processor_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|b_non_empty~q ),
	.r_val(\r_val~0_combout ),
	.clk_clk(clk_clk));

processor_processor_jtag_uart_scfifo_r the_processor_jtag_uart_scfifo_r(
	.q_b_0(q_b_0),
	.q_b_5(q_b_5),
	.q_b_4(q_b_4),
	.q_b_6(q_b_6),
	.q_b_7(q_b_7),
	.q_b_3(q_b_3),
	.q_b_2(q_b_2),
	.q_b_1(q_b_1),
	.r_sync_rst(r_sync_rst),
	.b_full(b_full),
	.counter_reg_bit_0(counter_reg_bit_0),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_4(counter_reg_bit_4),
	.b_non_empty(b_non_empty),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_1(counter_reg_bit_1),
	.fifo_rd(\fifo_rd~2_combout ),
	.t_ena(\processor_jtag_uart_alt_jtag_atlantic|t_ena~q ),
	.wr_rfifo(\wr_rfifo~combout ),
	.wdata_0(\processor_jtag_uart_alt_jtag_atlantic|wdata[0]~q ),
	.wdata_5(\processor_jtag_uart_alt_jtag_atlantic|wdata[5]~q ),
	.wdata_4(\processor_jtag_uart_alt_jtag_atlantic|wdata[4]~q ),
	.wdata_6(\processor_jtag_uart_alt_jtag_atlantic|wdata[6]~q ),
	.wdata_7(\processor_jtag_uart_alt_jtag_atlantic|wdata[7]~q ),
	.wdata_3(\processor_jtag_uart_alt_jtag_atlantic|wdata[3]~q ),
	.wdata_2(\processor_jtag_uart_alt_jtag_atlantic|wdata[2]~q ),
	.wdata_1(\processor_jtag_uart_alt_jtag_atlantic|wdata[1]~q ),
	.clk_clk(clk_clk));

processor_alt_jtag_atlantic processor_jtag_uart_alt_jtag_atlantic(
	.r_dat({\the_processor_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[7] ,\the_processor_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[6] ,\the_processor_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[5] ,
\the_processor_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[4] ,\the_processor_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[3] ,\the_processor_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[2] ,
\the_processor_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[1] ,\the_processor_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|FIFOram|q_b[0] }),
	.tdo1(tdo),
	.rst_n(r_sync_rst),
	.clr_break_line(clr_break_line),
	.t_dav(\t_dav~q ),
	.r_val(\r_val~q ),
	.t_pause1(\processor_jtag_uart_alt_jtag_atlantic|t_pause~q ),
	.rvalid01(\processor_jtag_uart_alt_jtag_atlantic|rvalid0~1_combout ),
	.t_ena1(\processor_jtag_uart_alt_jtag_atlantic|t_ena~q ),
	.wdata_0(\processor_jtag_uart_alt_jtag_atlantic|wdata[0]~q ),
	.wdata_5(\processor_jtag_uart_alt_jtag_atlantic|wdata[5]~q ),
	.wdata_4(\processor_jtag_uart_alt_jtag_atlantic|wdata[4]~q ),
	.wdata_6(\processor_jtag_uart_alt_jtag_atlantic|wdata[6]~q ),
	.wdata_7(\processor_jtag_uart_alt_jtag_atlantic|wdata[7]~q ),
	.wdata_3(\processor_jtag_uart_alt_jtag_atlantic|wdata[3]~q ),
	.wdata_2(\processor_jtag_uart_alt_jtag_atlantic|wdata[2]~q ),
	.wdata_1(\processor_jtag_uart_alt_jtag_atlantic|wdata[1]~q ),
	.altera_internal_jtag(altera_internal_jtag),
	.altera_internal_jtag1(altera_internal_jtag1),
	.state_4(state_4),
	.splitter_nodes_receive_0_3(splitter_nodes_receive_0_3),
	.virtual_ir_scan_reg(virtual_ir_scan_reg),
	.clr_reg(clr_reg),
	.state_3(state_3),
	.state_8(state_8),
	.irf_reg_0_1(irf_reg_0_1),
	.clk(clk_clk));

dffeas t_dav(
	.clk(clk_clk),
	.d(b_full),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\t_dav~q ),
	.prn(vcc));
defparam t_dav.is_wysiwyg = "true";
defparam t_dav.power_up = "low";

dffeas r_val(
	.clk(clk_clk),
	.d(\r_val~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\r_val~q ),
	.prn(vcc));
defparam r_val.is_wysiwyg = "true";
defparam r_val.power_up = "low";

dffeas fifo_wr(
	.clk(clk_clk),
	.d(\fifo_wr~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\fifo_wr~q ),
	.prn(vcc));
defparam fifo_wr.is_wysiwyg = "true";
defparam fifo_wr.power_up = "low";

cyclonev_lcell_comb \r_val~0 (
	.dataa(!\processor_jtag_uart_alt_jtag_atlantic|rvalid0~1_combout ),
	.datab(!\the_processor_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|b_non_empty~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\r_val~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \r_val~0 .extended_lut = "off";
defparam \r_val~0 .lut_mask = 64'h7777777777777777;
defparam \r_val~0 .shared_arith = "off";

cyclonev_lcell_comb \fifo_rd~2 (
	.dataa(!b_non_empty),
	.datab(!\fifo_rd~1_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fifo_rd~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fifo_rd~2 .extended_lut = "off";
defparam \fifo_rd~2 .lut_mask = 64'h7777777777777777;
defparam \fifo_rd~2 .shared_arith = "off";

cyclonev_lcell_comb wr_rfifo(
	.dataa(!b_full),
	.datab(!\processor_jtag_uart_alt_jtag_atlantic|t_ena~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wr_rfifo~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam wr_rfifo.extended_lut = "off";
defparam wr_rfifo.lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam wr_rfifo.shared_arith = "off";

cyclonev_lcell_comb \fifo_wr~0 (
	.dataa(!M_alu_result_2),
	.datab(!d_write),
	.datac(!\av_waitrequest~0_combout ),
	.datad(!b_full1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fifo_wr~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fifo_wr~0 .extended_lut = "off";
defparam \fifo_wr~0 .lut_mask = 64'hFFBFFFBFFFBFFFBF;
defparam \fifo_wr~0 .shared_arith = "off";

cyclonev_lcell_comb \Add1~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\the_processor_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Add1),
	.cout(\Add1~2 ),
	.shareout());
defparam \Add1~1 .extended_lut = "off";
defparam \Add1~1 .lut_mask = 64'h000000000000FF00;
defparam \Add1~1 .shared_arith = "off";

cyclonev_lcell_comb \Add1~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\the_processor_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(Add11),
	.cout(\Add1~6 ),
	.shareout());
defparam \Add1~5 .extended_lut = "off";
defparam \Add1~5 .lut_mask = 64'h000000000000FF00;
defparam \Add1~5 .shared_arith = "off";

cyclonev_lcell_comb \Add1~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\the_processor_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(Add12),
	.cout(\Add1~10 ),
	.shareout());
defparam \Add1~9 .extended_lut = "off";
defparam \Add1~9 .lut_mask = 64'h000000000000FF00;
defparam \Add1~9 .shared_arith = "off";

cyclonev_lcell_comb \Add1~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!b_full1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(Add13),
	.cout(),
	.shareout());
defparam \Add1~13 .extended_lut = "off";
defparam \Add1~13 .lut_mask = 64'h000000000000FF00;
defparam \Add1~13 .shared_arith = "off";

cyclonev_lcell_comb \Add1~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\the_processor_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(Add14),
	.cout(\Add1~18 ),
	.shareout());
defparam \Add1~17 .extended_lut = "off";
defparam \Add1~17 .lut_mask = 64'h000000000000FF00;
defparam \Add1~17 .shared_arith = "off";

cyclonev_lcell_comb \Add1~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\the_processor_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(Add15),
	.cout(\Add1~22 ),
	.shareout());
defparam \Add1~21 .extended_lut = "off";
defparam \Add1~21 .lut_mask = 64'h000000000000FF00;
defparam \Add1~21 .shared_arith = "off";

cyclonev_lcell_comb \Add1~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\the_processor_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(Add16),
	.cout(\Add1~26 ),
	.shareout());
defparam \Add1~25 .extended_lut = "off";
defparam \Add1~25 .lut_mask = 64'h000000000000FF00;
defparam \Add1~25 .shared_arith = "off";

dffeas av_waitrequest(
	.clk(clk_clk),
	.d(\av_waitrequest~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_waitrequest1),
	.prn(vcc));
defparam av_waitrequest.is_wysiwyg = "true";
defparam av_waitrequest.power_up = "low";

dffeas ien_AE(
	.clk(clk_clk),
	.d(M_st_data_1),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ien_AE~0_combout ),
	.q(ien_AE1),
	.prn(vcc));
defparam ien_AE.is_wysiwyg = "true";
defparam ien_AE.power_up = "low";

cyclonev_lcell_comb \av_readdata[9] (
	.dataa(!\fifo_AE~q ),
	.datab(!ien_AE1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(av_readdata_9),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_readdata[9] .extended_lut = "off";
defparam \av_readdata[9] .lut_mask = 64'h7777777777777777;
defparam \av_readdata[9] .shared_arith = "off";

dffeas ien_AF(
	.clk(clk_clk),
	.d(M_st_data_0),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ien_AE~0_combout ),
	.q(ien_AF1),
	.prn(vcc));
defparam ien_AF.is_wysiwyg = "true";
defparam ien_AF.power_up = "low";

cyclonev_lcell_comb \av_readdata[8]~0 (
	.dataa(!ien_AF1),
	.datab(!\pause_irq~q ),
	.datac(!\fifo_AF~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(av_readdata_8),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_readdata[8]~0 .extended_lut = "off";
defparam \av_readdata[8]~0 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \av_readdata[8]~0 .shared_arith = "off";

dffeas read_0(
	.clk(clk_clk),
	.d(\fifo_rd~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_01),
	.prn(vcc));
defparam read_0.is_wysiwyg = "true";
defparam read_0.power_up = "low";

dffeas woverflow(
	.clk(clk_clk),
	.d(\woverflow~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(woverflow1),
	.prn(vcc));
defparam woverflow.is_wysiwyg = "true";
defparam woverflow.power_up = "low";

dffeas rvalid(
	.clk(clk_clk),
	.d(\rvalid~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(rvalid1),
	.prn(vcc));
defparam rvalid.is_wysiwyg = "true";
defparam rvalid.power_up = "low";

dffeas ac(
	.clk(clk_clk),
	.d(\ac~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(ac1),
	.prn(vcc));
defparam ac.is_wysiwyg = "true";
defparam ac.power_up = "low";

cyclonev_lcell_comb \av_waitrequest~0 (
	.dataa(!Equal1),
	.datab(!Equal2),
	.datac(!av_waitrequest1),
	.datad(!Equal6),
	.datae(!read_latency_shift_reg),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_waitrequest~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_waitrequest~0 .extended_lut = "off";
defparam \av_waitrequest~0 .lut_mask = 64'hF7FFFFFFF7FFFFFF;
defparam \av_waitrequest~0 .shared_arith = "off";

cyclonev_lcell_comb \av_waitrequest~1 (
	.dataa(!d_write),
	.datab(!uav_read),
	.datac(!\av_waitrequest~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_waitrequest~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_waitrequest~1 .extended_lut = "off";
defparam \av_waitrequest~1 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \av_waitrequest~1 .shared_arith = "off";

cyclonev_lcell_comb \ien_AE~0 (
	.dataa(!M_alu_result_2),
	.datab(!d_write),
	.datac(!\av_waitrequest~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ien_AE~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ien_AE~0 .extended_lut = "off";
defparam \ien_AE~0 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \ien_AE~0 .shared_arith = "off";

cyclonev_lcell_comb \LessThan0~0 (
	.dataa(!\the_processor_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[0]~q ),
	.datab(!\the_processor_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[3]~q ),
	.datac(!\the_processor_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[2]~q ),
	.datad(!\the_processor_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan0~0 .extended_lut = "off";
defparam \LessThan0~0 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \LessThan0~0 .shared_arith = "off";

cyclonev_lcell_comb \LessThan0~1 (
	.dataa(!\the_processor_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[5]~q ),
	.datab(!\the_processor_jtag_uart_scfifo_w|wfifo|auto_generated|dpfifo|fifo_state|count_usedw|counter_reg_bit[4]~q ),
	.datac(!b_full1),
	.datad(!\LessThan0~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan0~1 .extended_lut = "off";
defparam \LessThan0~1 .lut_mask = 64'hFFFEFFFEFFFEFFFE;
defparam \LessThan0~1 .shared_arith = "off";

dffeas fifo_AE(
	.clk(clk_clk),
	.d(\LessThan0~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\fifo_AE~q ),
	.prn(vcc));
defparam fifo_AE.is_wysiwyg = "true";
defparam fifo_AE.power_up = "low";

cyclonev_lcell_comb \pause_irq~0 (
	.dataa(!\pause_irq~q ),
	.datab(!read_01),
	.datac(!b_non_empty),
	.datad(!\processor_jtag_uart_alt_jtag_atlantic|t_pause~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pause_irq~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pause_irq~0 .extended_lut = "off";
defparam \pause_irq~0 .lut_mask = 64'hDFFFDFFFDFFFDFFF;
defparam \pause_irq~0 .shared_arith = "off";

dffeas pause_irq(
	.clk(clk_clk),
	.d(\pause_irq~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\pause_irq~q ),
	.prn(vcc));
defparam pause_irq.is_wysiwyg = "true";
defparam pause_irq.power_up = "low";

cyclonev_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_0),
	.datae(gnd),
	.dataf(!counter_reg_bit_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout());
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~21 .shared_arith = "off";

cyclonev_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout());
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h000000000000FF00;
defparam \Add0~25 .shared_arith = "off";

cyclonev_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout());
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h000000000000FF00;
defparam \Add0~17 .shared_arith = "off";

cyclonev_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_4),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(\Add0~2 ),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h000000000000FF00;
defparam \Add0~1 .shared_arith = "off";

cyclonev_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_5),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout());
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h000000000000FF00;
defparam \Add0~5 .shared_arith = "off";

cyclonev_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!b_full),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout());
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h000000000000FF00;
defparam \Add0~9 .shared_arith = "off";

cyclonev_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(),
	.shareout());
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h0000000000000000;
defparam \Add0~13 .shared_arith = "off";

cyclonev_lcell_comb \LessThan1~0 (
	.dataa(!counter_reg_bit_0),
	.datab(!\Add0~17_sumout ),
	.datac(!\Add0~21_sumout ),
	.datad(!\Add0~25_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan1~0 .extended_lut = "off";
defparam \LessThan1~0 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \LessThan1~0 .shared_arith = "off";

cyclonev_lcell_comb \LessThan1~1 (
	.dataa(!\Add0~1_sumout ),
	.datab(!\Add0~5_sumout ),
	.datac(!\Add0~9_sumout ),
	.datad(!\Add0~13_sumout ),
	.datae(!\LessThan1~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan1~1 .extended_lut = "off";
defparam \LessThan1~1 .lut_mask = 64'hFFFFFFFEFFFFFFFE;
defparam \LessThan1~1 .shared_arith = "off";

dffeas fifo_AF(
	.clk(clk_clk),
	.d(\LessThan1~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\fifo_AF~q ),
	.prn(vcc));
defparam fifo_AF.is_wysiwyg = "true";
defparam fifo_AF.power_up = "low";

cyclonev_lcell_comb \fifo_rd~0 (
	.dataa(!M_alu_result_2),
	.datab(!d_read),
	.datac(!read_accepted),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fifo_rd~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fifo_rd~0 .extended_lut = "off";
defparam \fifo_rd~0 .lut_mask = 64'hFBFBFBFBFBFBFBFB;
defparam \fifo_rd~0 .shared_arith = "off";

cyclonev_lcell_comb \fifo_rd~1 (
	.dataa(!Equal1),
	.datab(!Equal2),
	.datac(!av_waitrequest1),
	.datad(!Equal6),
	.datae(!read_latency_shift_reg),
	.dataf(!\fifo_rd~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\fifo_rd~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \fifo_rd~1 .extended_lut = "off";
defparam \fifo_rd~1 .lut_mask = 64'hF7FFFFFFFFFFFFFF;
defparam \fifo_rd~1 .shared_arith = "off";

cyclonev_lcell_comb \woverflow~0 (
	.dataa(!M_alu_result_2),
	.datab(!d_write),
	.datac(!\av_waitrequest~0_combout ),
	.datad(!b_full1),
	.datae(!woverflow1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\woverflow~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \woverflow~0 .extended_lut = "off";
defparam \woverflow~0 .lut_mask = 64'h96FFFFFF96FFFFFF;
defparam \woverflow~0 .shared_arith = "off";

cyclonev_lcell_comb \rvalid~0 (
	.dataa(!b_non_empty),
	.datab(!rvalid1),
	.datac(!\fifo_rd~1_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rvalid~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rvalid~0 .extended_lut = "off";
defparam \rvalid~0 .lut_mask = 64'h5353535353535353;
defparam \rvalid~0 .shared_arith = "off";

cyclonev_lcell_comb \ac~0 (
	.dataa(!ac1),
	.datab(!M_st_data_10),
	.datac(!\ien_AE~0_combout ),
	.datad(!\processor_jtag_uart_alt_jtag_atlantic|t_pause~q ),
	.datae(!\processor_jtag_uart_alt_jtag_atlantic|t_ena~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ac~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ac~0 .extended_lut = "off";
defparam \ac~0 .lut_mask = 64'hFDFFFFFFFDFFFFFF;
defparam \ac~0 .shared_arith = "off";

endmodule

module processor_alt_jtag_atlantic (
	r_dat,
	tdo1,
	rst_n,
	clr_break_line,
	t_dav,
	r_val,
	t_pause1,
	rvalid01,
	t_ena1,
	wdata_0,
	wdata_5,
	wdata_4,
	wdata_6,
	wdata_7,
	wdata_3,
	wdata_2,
	wdata_1,
	altera_internal_jtag,
	altera_internal_jtag1,
	state_4,
	splitter_nodes_receive_0_3,
	virtual_ir_scan_reg,
	clr_reg,
	state_3,
	state_8,
	irf_reg_0_1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	[7:0] r_dat;
output 	tdo1;
input 	rst_n;
input 	clr_break_line;
input 	t_dav;
input 	r_val;
output 	t_pause1;
output 	rvalid01;
output 	t_ena1;
output 	wdata_0;
output 	wdata_5;
output 	wdata_4;
output 	wdata_6;
output 	wdata_7;
output 	wdata_3;
output 	wdata_2;
output 	wdata_1;
input 	altera_internal_jtag;
input 	altera_internal_jtag1;
input 	state_4;
input 	splitter_nodes_receive_0_3;
input 	virtual_ir_scan_reg;
input 	clr_reg;
input 	state_3;
input 	state_8;
input 	irf_reg_0_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \state~1_combout ;
wire \state~q ;
wire \td_shift[0]~2_combout ;
wire \count[2]~q ;
wire \count[3]~q ;
wire \count[4]~q ;
wire \count[5]~q ;
wire \count[6]~q ;
wire \count[7]~q ;
wire \count[8]~q ;
wire \count[9]~0_combout ;
wire \count[9]~q ;
wire \count[9]~_wirecell_combout ;
wire \count[0]~q ;
wire \count[1]~q ;
wire \state~0_combout ;
wire \user_saw_rvalid~0_combout ;
wire \user_saw_rvalid~q ;
wire \td_shift[10]~q ;
wire \r_ena1~q ;
wire \r_ena~0_combout ;
wire \rdata[7]~q ;
wire \td_shift~3_combout ;
wire \td_shift[9]~q ;
wire \td_shift~0_combout ;
wire \tck_t_dav~0_combout ;
wire \tck_t_dav~q ;
wire \write_stalled~0_combout ;
wire \write_stalled~1_combout ;
wire \write_stalled~q ;
wire \td_shift~4_combout ;
wire \rdata[0]~q ;
wire \rdata[6]~q ;
wire \td_shift~10_combout ;
wire \td_shift[8]~q ;
wire \rdata[5]~q ;
wire \td_shift~11_combout ;
wire \td_shift[7]~q ;
wire \rdata[4]~q ;
wire \td_shift~12_combout ;
wire \td_shift[6]~q ;
wire \rdata[3]~q ;
wire \td_shift~9_combout ;
wire \td_shift[5]~q ;
wire \rdata[2]~q ;
wire \td_shift~8_combout ;
wire \td_shift[4]~q ;
wire \rdata[1]~q ;
wire \td_shift~7_combout ;
wire \td_shift[3]~q ;
wire \td_shift~6_combout ;
wire \td_shift[2]~q ;
wire \td_shift~5_combout ;
wire \td_shift[1]~q ;
wire \read_req~q ;
wire \read~0_combout ;
wire \read~q ;
wire \read1~q ;
wire \read2~q ;
wire \always2~0_combout ;
wire \rst2~q ;
wire \rvalid0~0_combout ;
wire \rvalid0~q ;
wire \rvalid~q ;
wire \td_shift~1_combout ;
wire \td_shift[0]~q ;
wire \jupdate~0_combout ;
wire \jupdate~q ;
wire \jupdate1~q ;
wire \jupdate2~q ;
wire \always2~1_combout ;
wire \write~0_combout ;
wire \wdata[7]~0_combout ;
wire \write~q ;
wire \write1~q ;
wire \write2~q ;
wire \always2~2_combout ;
wire \write_valid~q ;
wire \t_pause~0_combout ;
wire \t_ena~0_combout ;


dffeas tdo(
	.clk(!altera_internal_jtag),
	.d(\td_shift[0]~q ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(tdo1),
	.prn(vcc));
defparam tdo.is_wysiwyg = "true";
defparam tdo.power_up = "low";

dffeas t_pause(
	.clk(clk),
	.d(\t_pause~0_combout ),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(t_pause1),
	.prn(vcc));
defparam t_pause.is_wysiwyg = "true";
defparam t_pause.power_up = "low";

cyclonev_lcell_comb \rvalid0~1 (
	.dataa(!\rvalid0~q ),
	.datab(!\r_ena~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(rvalid01),
	.sumout(),
	.cout(),
	.shareout());
defparam \rvalid0~1 .extended_lut = "off";
defparam \rvalid0~1 .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \rvalid0~1 .shared_arith = "off";

dffeas t_ena(
	.clk(clk),
	.d(\t_ena~0_combout ),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(t_ena1),
	.prn(vcc));
defparam t_ena.is_wysiwyg = "true";
defparam t_ena.power_up = "low";

dffeas \wdata[0] (
	.clk(altera_internal_jtag),
	.d(altera_internal_jtag1),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_stalled~1_combout ),
	.q(wdata_0),
	.prn(vcc));
defparam \wdata[0] .is_wysiwyg = "true";
defparam \wdata[0] .power_up = "low";

dffeas \wdata[5] (
	.clk(altera_internal_jtag),
	.d(\td_shift[9]~q ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wdata[7]~0_combout ),
	.q(wdata_5),
	.prn(vcc));
defparam \wdata[5] .is_wysiwyg = "true";
defparam \wdata[5] .power_up = "low";

dffeas \wdata[4] (
	.clk(altera_internal_jtag),
	.d(\td_shift[8]~q ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wdata[7]~0_combout ),
	.q(wdata_4),
	.prn(vcc));
defparam \wdata[4] .is_wysiwyg = "true";
defparam \wdata[4] .power_up = "low";

dffeas \wdata[6] (
	.clk(altera_internal_jtag),
	.d(\td_shift[10]~q ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wdata[7]~0_combout ),
	.q(wdata_6),
	.prn(vcc));
defparam \wdata[6] .is_wysiwyg = "true";
defparam \wdata[6] .power_up = "low";

dffeas \wdata[7] (
	.clk(altera_internal_jtag),
	.d(altera_internal_jtag1),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wdata[7]~0_combout ),
	.q(wdata_7),
	.prn(vcc));
defparam \wdata[7] .is_wysiwyg = "true";
defparam \wdata[7] .power_up = "low";

dffeas \wdata[3] (
	.clk(altera_internal_jtag),
	.d(\td_shift[7]~q ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wdata[7]~0_combout ),
	.q(wdata_3),
	.prn(vcc));
defparam \wdata[3] .is_wysiwyg = "true";
defparam \wdata[3] .power_up = "low";

dffeas \wdata[2] (
	.clk(altera_internal_jtag),
	.d(\td_shift[6]~q ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wdata[7]~0_combout ),
	.q(wdata_2),
	.prn(vcc));
defparam \wdata[2] .is_wysiwyg = "true";
defparam \wdata[2] .power_up = "low";

dffeas \wdata[1] (
	.clk(altera_internal_jtag),
	.d(\td_shift[5]~q ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wdata[7]~0_combout ),
	.q(wdata_1),
	.prn(vcc));
defparam \wdata[1] .is_wysiwyg = "true";
defparam \wdata[1] .power_up = "low";

cyclonev_lcell_comb \state~1 (
	.dataa(!virtual_ir_scan_reg),
	.datab(!splitter_nodes_receive_0_3),
	.datac(!state_3),
	.datad(!state_4),
	.datae(!\state~q ),
	.dataf(!altera_internal_jtag1),
	.datag(!irf_reg_0_1),
	.cin(gnd),
	.sharein(gnd),
	.combout(\state~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \state~1 .extended_lut = "on";
defparam \state~1 .lut_mask = 64'hFF6FFF6FFF6FFF6F;
defparam \state~1 .shared_arith = "off";

dffeas state(
	.clk(altera_internal_jtag),
	.d(\state~1_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state~q ),
	.prn(vcc));
defparam state.is_wysiwyg = "true";
defparam state.power_up = "low";

cyclonev_lcell_comb \td_shift[0]~2 (
	.dataa(!state_4),
	.datab(!splitter_nodes_receive_0_3),
	.datac(!virtual_ir_scan_reg),
	.datad(!state_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\td_shift[0]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \td_shift[0]~2 .extended_lut = "off";
defparam \td_shift[0]~2 .lut_mask = 64'hF7FFF7FFF7FFF7FF;
defparam \td_shift[0]~2 .shared_arith = "off";

dffeas \count[2] (
	.clk(altera_internal_jtag),
	.d(\count[1]~q ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(!state_4),
	.sload(gnd),
	.ena(\td_shift[0]~2_combout ),
	.q(\count[2]~q ),
	.prn(vcc));
defparam \count[2] .is_wysiwyg = "true";
defparam \count[2] .power_up = "low";

dffeas \count[3] (
	.clk(altera_internal_jtag),
	.d(\count[2]~q ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(!state_4),
	.sload(gnd),
	.ena(\td_shift[0]~2_combout ),
	.q(\count[3]~q ),
	.prn(vcc));
defparam \count[3] .is_wysiwyg = "true";
defparam \count[3] .power_up = "low";

dffeas \count[4] (
	.clk(altera_internal_jtag),
	.d(\count[3]~q ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(!state_4),
	.sload(gnd),
	.ena(\td_shift[0]~2_combout ),
	.q(\count[4]~q ),
	.prn(vcc));
defparam \count[4] .is_wysiwyg = "true";
defparam \count[4] .power_up = "low";

dffeas \count[5] (
	.clk(altera_internal_jtag),
	.d(\count[4]~q ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(!state_4),
	.sload(gnd),
	.ena(\td_shift[0]~2_combout ),
	.q(\count[5]~q ),
	.prn(vcc));
defparam \count[5] .is_wysiwyg = "true";
defparam \count[5] .power_up = "low";

dffeas \count[6] (
	.clk(altera_internal_jtag),
	.d(\count[5]~q ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(!state_4),
	.sload(gnd),
	.ena(\td_shift[0]~2_combout ),
	.q(\count[6]~q ),
	.prn(vcc));
defparam \count[6] .is_wysiwyg = "true";
defparam \count[6] .power_up = "low";

dffeas \count[7] (
	.clk(altera_internal_jtag),
	.d(\count[6]~q ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(!state_4),
	.sload(gnd),
	.ena(\td_shift[0]~2_combout ),
	.q(\count[7]~q ),
	.prn(vcc));
defparam \count[7] .is_wysiwyg = "true";
defparam \count[7] .power_up = "low";

dffeas \count[8] (
	.clk(altera_internal_jtag),
	.d(\count[7]~q ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(!state_4),
	.sload(gnd),
	.ena(\td_shift[0]~2_combout ),
	.q(\count[8]~q ),
	.prn(vcc));
defparam \count[8] .is_wysiwyg = "true";
defparam \count[8] .power_up = "low";

cyclonev_lcell_comb \count[9]~0 (
	.dataa(!irf_reg_0_1),
	.datab(!\state~q ),
	.datac(!altera_internal_jtag1),
	.datad(!state_4),
	.datae(!\count[8]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\count[9]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \count[9]~0 .extended_lut = "off";
defparam \count[9]~0 .lut_mask = 64'hFFFFFFF7FFFFFFF7;
defparam \count[9]~0 .shared_arith = "off";

dffeas \count[9] (
	.clk(altera_internal_jtag),
	.d(\count[9]~0_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\td_shift[0]~2_combout ),
	.q(\count[9]~q ),
	.prn(vcc));
defparam \count[9] .is_wysiwyg = "true";
defparam \count[9] .power_up = "low";

cyclonev_lcell_comb \count[9]~_wirecell (
	.dataa(!\count[9]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\count[9]~_wirecell_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \count[9]~_wirecell .extended_lut = "off";
defparam \count[9]~_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \count[9]~_wirecell .shared_arith = "off";

dffeas \count[0] (
	.clk(altera_internal_jtag),
	.d(\count[9]~_wirecell_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(!state_4),
	.sload(gnd),
	.ena(\td_shift[0]~2_combout ),
	.q(\count[0]~q ),
	.prn(vcc));
defparam \count[0] .is_wysiwyg = "true";
defparam \count[0] .power_up = "low";

dffeas \count[1] (
	.clk(altera_internal_jtag),
	.d(\count[0]~q ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(!state_4),
	.sload(gnd),
	.ena(\td_shift[0]~2_combout ),
	.q(\count[1]~q ),
	.prn(vcc));
defparam \count[1] .is_wysiwyg = "true";
defparam \count[1] .power_up = "low";

cyclonev_lcell_comb \state~0 (
	.dataa(!state_4),
	.datab(!splitter_nodes_receive_0_3),
	.datac(!virtual_ir_scan_reg),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\state~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \state~0 .extended_lut = "off";
defparam \state~0 .lut_mask = 64'hF7F7F7F7F7F7F7F7;
defparam \state~0 .shared_arith = "off";

cyclonev_lcell_comb \user_saw_rvalid~0 (
	.dataa(!irf_reg_0_1),
	.datab(!\td_shift[0]~q ),
	.datac(!\state~q ),
	.datad(!\user_saw_rvalid~q ),
	.datae(!\state~0_combout ),
	.dataf(!\count[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\user_saw_rvalid~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \user_saw_rvalid~0 .extended_lut = "off";
defparam \user_saw_rvalid~0 .lut_mask = 64'h7BFFB7FFB7FF7BFF;
defparam \user_saw_rvalid~0 .shared_arith = "off";

dffeas user_saw_rvalid(
	.clk(altera_internal_jtag),
	.d(\user_saw_rvalid~0_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\user_saw_rvalid~q ),
	.prn(vcc));
defparam user_saw_rvalid.is_wysiwyg = "true";
defparam user_saw_rvalid.power_up = "low";

dffeas \td_shift[10] (
	.clk(altera_internal_jtag),
	.d(altera_internal_jtag1),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(!state_4),
	.sload(gnd),
	.ena(\td_shift[0]~2_combout ),
	.q(\td_shift[10]~q ),
	.prn(vcc));
defparam \td_shift[10] .is_wysiwyg = "true";
defparam \td_shift[10] .power_up = "low";

dffeas r_ena1(
	.clk(clk),
	.d(rvalid01),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\r_ena1~q ),
	.prn(vcc));
defparam r_ena1.is_wysiwyg = "true";
defparam r_ena1.power_up = "low";

cyclonev_lcell_comb \r_ena~0 (
	.dataa(!r_val),
	.datab(!\r_ena1~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\r_ena~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \r_ena~0 .extended_lut = "off";
defparam \r_ena~0 .lut_mask = 64'h7777777777777777;
defparam \r_ena~0 .shared_arith = "off";

dffeas \rdata[7] (
	.clk(clk),
	.d(r_dat[7]),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\r_ena~0_combout ),
	.q(\rdata[7]~q ),
	.prn(vcc));
defparam \rdata[7] .is_wysiwyg = "true";
defparam \rdata[7] .power_up = "low";

cyclonev_lcell_comb \td_shift~3 (
	.dataa(!\count[9]~q ),
	.datab(!\td_shift[10]~q ),
	.datac(!\rdata[7]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\td_shift~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \td_shift~3 .extended_lut = "off";
defparam \td_shift~3 .lut_mask = 64'h2727272727272727;
defparam \td_shift~3 .shared_arith = "off";

dffeas \td_shift[9] (
	.clk(altera_internal_jtag),
	.d(\td_shift~3_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(!state_4),
	.sload(gnd),
	.ena(\td_shift[0]~2_combout ),
	.q(\td_shift[9]~q ),
	.prn(vcc));
defparam \td_shift[9] .is_wysiwyg = "true";
defparam \td_shift[9] .power_up = "low";

cyclonev_lcell_comb \td_shift~0 (
	.dataa(!irf_reg_0_1),
	.datab(!\state~q ),
	.datac(!\count[1]~q ),
	.datad(!\user_saw_rvalid~q ),
	.datae(!\td_shift[9]~q ),
	.dataf(!altera_internal_jtag1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\td_shift~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \td_shift~0 .extended_lut = "off";
defparam \td_shift~0 .lut_mask = 64'hFFFFBF8FFFFFFFFF;
defparam \td_shift~0 .shared_arith = "off";

cyclonev_lcell_comb \tck_t_dav~0 (
	.dataa(!t_dav),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\tck_t_dav~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \tck_t_dav~0 .extended_lut = "off";
defparam \tck_t_dav~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \tck_t_dav~0 .shared_arith = "off";

dffeas tck_t_dav(
	.clk(altera_internal_jtag),
	.d(\tck_t_dav~0_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\tck_t_dav~q ),
	.prn(vcc));
defparam tck_t_dav.is_wysiwyg = "true";
defparam tck_t_dav.power_up = "low";

cyclonev_lcell_comb \write_stalled~0 (
	.dataa(!altera_internal_jtag1),
	.datab(!\tck_t_dav~q ),
	.datac(!\td_shift[10]~q ),
	.datad(!\write_stalled~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\write_stalled~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \write_stalled~0 .extended_lut = "off";
defparam \write_stalled~0 .lut_mask = 64'hEFFFEFFFEFFFEFFF;
defparam \write_stalled~0 .shared_arith = "off";

cyclonev_lcell_comb \write_stalled~1 (
	.dataa(!irf_reg_0_1),
	.datab(!\state~q ),
	.datac(!\count[1]~q ),
	.datad(!state_4),
	.datae(!splitter_nodes_receive_0_3),
	.dataf(!virtual_ir_scan_reg),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\write_stalled~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \write_stalled~1 .extended_lut = "off";
defparam \write_stalled~1 .lut_mask = 64'hFFFFFFFFBFFFFFFF;
defparam \write_stalled~1 .shared_arith = "off";

dffeas write_stalled(
	.clk(altera_internal_jtag),
	.d(\write_stalled~0_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_stalled~1_combout ),
	.q(\write_stalled~q ),
	.prn(vcc));
defparam write_stalled.is_wysiwyg = "true";
defparam write_stalled.power_up = "low";

cyclonev_lcell_comb \td_shift~4 (
	.dataa(!irf_reg_0_1),
	.datab(!\state~q ),
	.datac(!\count[1]~q ),
	.datad(!\user_saw_rvalid~q ),
	.datae(!\td_shift[9]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\td_shift~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \td_shift~4 .extended_lut = "off";
defparam \td_shift~4 .lut_mask = 64'hFFFFFFBFFFFFFFBF;
defparam \td_shift~4 .shared_arith = "off";

dffeas \rdata[0] (
	.clk(clk),
	.d(r_dat[0]),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\r_ena~0_combout ),
	.q(\rdata[0]~q ),
	.prn(vcc));
defparam \rdata[0] .is_wysiwyg = "true";
defparam \rdata[0] .power_up = "low";

dffeas \rdata[6] (
	.clk(clk),
	.d(r_dat[6]),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\r_ena~0_combout ),
	.q(\rdata[6]~q ),
	.prn(vcc));
defparam \rdata[6] .is_wysiwyg = "true";
defparam \rdata[6] .power_up = "low";

cyclonev_lcell_comb \td_shift~10 (
	.dataa(!\td_shift[9]~q ),
	.datab(!\count[9]~q ),
	.datac(!\rdata[6]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\td_shift~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \td_shift~10 .extended_lut = "off";
defparam \td_shift~10 .lut_mask = 64'h4747474747474747;
defparam \td_shift~10 .shared_arith = "off";

dffeas \td_shift[8] (
	.clk(altera_internal_jtag),
	.d(\td_shift~10_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(!state_4),
	.sload(gnd),
	.ena(\td_shift[0]~2_combout ),
	.q(\td_shift[8]~q ),
	.prn(vcc));
defparam \td_shift[8] .is_wysiwyg = "true";
defparam \td_shift[8] .power_up = "low";

dffeas \rdata[5] (
	.clk(clk),
	.d(r_dat[5]),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\r_ena~0_combout ),
	.q(\rdata[5]~q ),
	.prn(vcc));
defparam \rdata[5] .is_wysiwyg = "true";
defparam \rdata[5] .power_up = "low";

cyclonev_lcell_comb \td_shift~11 (
	.dataa(!\count[9]~q ),
	.datab(!state_4),
	.datac(!\td_shift~4_combout ),
	.datad(!\td_shift[8]~q ),
	.datae(!\rdata[5]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\td_shift~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \td_shift~11 .extended_lut = "off";
defparam \td_shift~11 .lut_mask = 64'hB1FFFFFFB1FFFFFF;
defparam \td_shift~11 .shared_arith = "off";

dffeas \td_shift[7] (
	.clk(altera_internal_jtag),
	.d(\td_shift~11_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\td_shift[0]~2_combout ),
	.q(\td_shift[7]~q ),
	.prn(vcc));
defparam \td_shift[7] .is_wysiwyg = "true";
defparam \td_shift[7] .power_up = "low";

dffeas \rdata[4] (
	.clk(clk),
	.d(r_dat[4]),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\r_ena~0_combout ),
	.q(\rdata[4]~q ),
	.prn(vcc));
defparam \rdata[4] .is_wysiwyg = "true";
defparam \rdata[4] .power_up = "low";

cyclonev_lcell_comb \td_shift~12 (
	.dataa(!irf_reg_0_1),
	.datab(!\count[9]~q ),
	.datac(!state_4),
	.datad(!\td_shift~4_combout ),
	.datae(!\td_shift[7]~q ),
	.dataf(!\rdata[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\td_shift~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \td_shift~12 .extended_lut = "off";
defparam \td_shift~12 .lut_mask = 64'hFF7DFFFFFFFFFFFF;
defparam \td_shift~12 .shared_arith = "off";

dffeas \td_shift[6] (
	.clk(altera_internal_jtag),
	.d(\td_shift~12_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\td_shift[0]~2_combout ),
	.q(\td_shift[6]~q ),
	.prn(vcc));
defparam \td_shift[6] .is_wysiwyg = "true";
defparam \td_shift[6] .power_up = "low";

dffeas \rdata[3] (
	.clk(clk),
	.d(r_dat[3]),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\r_ena~0_combout ),
	.q(\rdata[3]~q ),
	.prn(vcc));
defparam \rdata[3] .is_wysiwyg = "true";
defparam \rdata[3] .power_up = "low";

cyclonev_lcell_comb \td_shift~9 (
	.dataa(!irf_reg_0_1),
	.datab(!\count[9]~q ),
	.datac(!state_4),
	.datad(!\td_shift~4_combout ),
	.datae(!\td_shift[6]~q ),
	.dataf(!\rdata[3]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\td_shift~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \td_shift~9 .extended_lut = "off";
defparam \td_shift~9 .lut_mask = 64'hFF7DFFFFFFFFFFFF;
defparam \td_shift~9 .shared_arith = "off";

dffeas \td_shift[5] (
	.clk(altera_internal_jtag),
	.d(\td_shift~9_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\td_shift[0]~2_combout ),
	.q(\td_shift[5]~q ),
	.prn(vcc));
defparam \td_shift[5] .is_wysiwyg = "true";
defparam \td_shift[5] .power_up = "low";

dffeas \rdata[2] (
	.clk(clk),
	.d(r_dat[2]),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\r_ena~0_combout ),
	.q(\rdata[2]~q ),
	.prn(vcc));
defparam \rdata[2] .is_wysiwyg = "true";
defparam \rdata[2] .power_up = "low";

cyclonev_lcell_comb \td_shift~8 (
	.dataa(!\count[9]~q ),
	.datab(!state_4),
	.datac(!\td_shift~4_combout ),
	.datad(!\td_shift[5]~q ),
	.datae(!\rdata[2]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\td_shift~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \td_shift~8 .extended_lut = "off";
defparam \td_shift~8 .lut_mask = 64'hB1FFFFFFB1FFFFFF;
defparam \td_shift~8 .shared_arith = "off";

dffeas \td_shift[4] (
	.clk(altera_internal_jtag),
	.d(\td_shift~8_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\td_shift[0]~2_combout ),
	.q(\td_shift[4]~q ),
	.prn(vcc));
defparam \td_shift[4] .is_wysiwyg = "true";
defparam \td_shift[4] .power_up = "low";

dffeas \rdata[1] (
	.clk(clk),
	.d(r_dat[1]),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\r_ena~0_combout ),
	.q(\rdata[1]~q ),
	.prn(vcc));
defparam \rdata[1] .is_wysiwyg = "true";
defparam \rdata[1] .power_up = "low";

cyclonev_lcell_comb \td_shift~7 (
	.dataa(!\count[9]~q ),
	.datab(!state_4),
	.datac(!\td_shift~4_combout ),
	.datad(!\td_shift[4]~q ),
	.datae(!\rdata[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\td_shift~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \td_shift~7 .extended_lut = "off";
defparam \td_shift~7 .lut_mask = 64'hB1FFFFFFB1FFFFFF;
defparam \td_shift~7 .shared_arith = "off";

dffeas \td_shift[3] (
	.clk(altera_internal_jtag),
	.d(\td_shift~7_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\td_shift[0]~2_combout ),
	.q(\td_shift[3]~q ),
	.prn(vcc));
defparam \td_shift[3] .is_wysiwyg = "true";
defparam \td_shift[3] .power_up = "low";

cyclonev_lcell_comb \td_shift~6 (
	.dataa(!irf_reg_0_1),
	.datab(!\count[9]~q ),
	.datac(!state_4),
	.datad(!\td_shift~4_combout ),
	.datae(!\rdata[0]~q ),
	.dataf(!\td_shift[3]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\td_shift~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \td_shift~6 .extended_lut = "off";
defparam \td_shift~6 .lut_mask = 64'hFF7DFFFFFFFFFFFF;
defparam \td_shift~6 .shared_arith = "off";

dffeas \td_shift[2] (
	.clk(altera_internal_jtag),
	.d(\td_shift~6_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\td_shift[0]~2_combout ),
	.q(\td_shift[2]~q ),
	.prn(vcc));
defparam \td_shift[2] .is_wysiwyg = "true";
defparam \td_shift[2] .power_up = "low";

cyclonev_lcell_comb \td_shift~5 (
	.dataa(!irf_reg_0_1),
	.datab(!\count[9]~q ),
	.datac(!state_4),
	.datad(!\write_stalled~q ),
	.datae(!\td_shift~4_combout ),
	.dataf(!\td_shift[2]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\td_shift~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \td_shift~5 .extended_lut = "off";
defparam \td_shift~5 .lut_mask = 64'hFFFF7DFFFFFFFFFF;
defparam \td_shift~5 .shared_arith = "off";

dffeas \td_shift[1] (
	.clk(altera_internal_jtag),
	.d(\td_shift~5_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\td_shift[0]~2_combout ),
	.q(\td_shift[1]~q ),
	.prn(vcc));
defparam \td_shift[1] .is_wysiwyg = "true";
defparam \td_shift[1] .power_up = "low";

dffeas read_req(
	.clk(altera_internal_jtag),
	.d(\td_shift[9]~q ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_stalled~1_combout ),
	.q(\read_req~q ),
	.prn(vcc));
defparam read_req.is_wysiwyg = "true";
defparam read_req.power_up = "low";

cyclonev_lcell_comb \read~0 (
	.dataa(!\read~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read~0 .extended_lut = "off";
defparam \read~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \read~0 .shared_arith = "off";

dffeas read(
	.clk(altera_internal_jtag),
	.d(\read~0_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_stalled~1_combout ),
	.q(\read~q ),
	.prn(vcc));
defparam read.is_wysiwyg = "true";
defparam read.power_up = "low";

dffeas read1(
	.clk(clk),
	.d(\read~q ),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\read1~q ),
	.prn(vcc));
defparam read1.is_wysiwyg = "true";
defparam read1.power_up = "low";

dffeas read2(
	.clk(clk),
	.d(\read1~q ),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\read2~q ),
	.prn(vcc));
defparam read2.is_wysiwyg = "true";
defparam read2.power_up = "low";

cyclonev_lcell_comb \always2~0 (
	.dataa(!\read1~q ),
	.datab(!\read2~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always2~0 .extended_lut = "off";
defparam \always2~0 .lut_mask = 64'h6666666666666666;
defparam \always2~0 .shared_arith = "off";

dffeas rst2(
	.clk(clk),
	.d(clr_break_line),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rst2~q ),
	.prn(vcc));
defparam rst2.is_wysiwyg = "true";
defparam rst2.power_up = "low";

cyclonev_lcell_comb \rvalid0~0 (
	.dataa(!\user_saw_rvalid~q ),
	.datab(!\rvalid0~q ),
	.datac(!\r_ena~0_combout ),
	.datad(!\read_req~q ),
	.datae(!\always2~0_combout ),
	.dataf(!\rst2~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rvalid0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rvalid0~0 .extended_lut = "off";
defparam \rvalid0~0 .lut_mask = 64'hFFFFFFFFFFFFFFBF;
defparam \rvalid0~0 .shared_arith = "off";

dffeas rvalid0(
	.clk(clk),
	.d(\rvalid0~0_combout ),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rvalid0~q ),
	.prn(vcc));
defparam rvalid0.is_wysiwyg = "true";
defparam rvalid0.power_up = "low";

dffeas rvalid(
	.clk(clk),
	.d(\rvalid0~q ),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rvalid~q ),
	.prn(vcc));
defparam rvalid.is_wysiwyg = "true";
defparam rvalid.power_up = "low";

cyclonev_lcell_comb \td_shift~1 (
	.dataa(!\state~q ),
	.datab(!\td_shift~0_combout ),
	.datac(!\tck_t_dav~q ),
	.datad(!\td_shift[1]~q ),
	.datae(!\count[9]~q ),
	.dataf(!\rvalid~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\td_shift~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \td_shift~1 .extended_lut = "off";
defparam \td_shift~1 .lut_mask = 64'hBFFFEFFFFFFFFFFF;
defparam \td_shift~1 .shared_arith = "off";

dffeas \td_shift[0] (
	.clk(altera_internal_jtag),
	.d(\td_shift~1_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(!state_4),
	.sload(gnd),
	.ena(\td_shift[0]~2_combout ),
	.q(\td_shift[0]~q ),
	.prn(vcc));
defparam \td_shift[0] .is_wysiwyg = "true";
defparam \td_shift[0] .power_up = "low";

cyclonev_lcell_comb \jupdate~0 (
	.dataa(!irf_reg_0_1),
	.datab(!splitter_nodes_receive_0_3),
	.datac(!virtual_ir_scan_reg),
	.datad(!\jupdate~q ),
	.datae(!state_8),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\jupdate~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \jupdate~0 .extended_lut = "off";
defparam \jupdate~0 .lut_mask = 64'h9669699696696996;
defparam \jupdate~0 .shared_arith = "off";

dffeas jupdate(
	.clk(!altera_internal_jtag),
	.d(\jupdate~0_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\jupdate~q ),
	.prn(vcc));
defparam jupdate.is_wysiwyg = "true";
defparam jupdate.power_up = "low";

dffeas jupdate1(
	.clk(clk),
	.d(\jupdate~q ),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\jupdate1~q ),
	.prn(vcc));
defparam jupdate1.is_wysiwyg = "true";
defparam jupdate1.power_up = "low";

dffeas jupdate2(
	.clk(clk),
	.d(\jupdate1~q ),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\jupdate2~q ),
	.prn(vcc));
defparam jupdate2.is_wysiwyg = "true";
defparam jupdate2.power_up = "low";

cyclonev_lcell_comb \always2~1 (
	.dataa(!\jupdate1~q ),
	.datab(!\jupdate2~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always2~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always2~1 .extended_lut = "off";
defparam \always2~1 .lut_mask = 64'h6666666666666666;
defparam \always2~1 .shared_arith = "off";

cyclonev_lcell_comb \write~0 (
	.dataa(!\write~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\write~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \write~0 .extended_lut = "off";
defparam \write~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \write~0 .shared_arith = "off";

cyclonev_lcell_comb \wdata[7]~0 (
	.dataa(!irf_reg_0_1),
	.datab(!\state~q ),
	.datac(!state_4),
	.datad(!splitter_nodes_receive_0_3),
	.datae(!virtual_ir_scan_reg),
	.dataf(!\count[8]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wdata[7]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wdata[7]~0 .extended_lut = "off";
defparam \wdata[7]~0 .lut_mask = 64'hFFFFBFFFFFFFFFFF;
defparam \wdata[7]~0 .shared_arith = "off";

dffeas write(
	.clk(altera_internal_jtag),
	.d(\write~0_combout ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\wdata[7]~0_combout ),
	.q(\write~q ),
	.prn(vcc));
defparam write.is_wysiwyg = "true";
defparam write.power_up = "low";

dffeas write1(
	.clk(clk),
	.d(\write~q ),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\write1~q ),
	.prn(vcc));
defparam write1.is_wysiwyg = "true";
defparam write1.power_up = "low";

dffeas write2(
	.clk(clk),
	.d(\write1~q ),
	.asdata(vcc),
	.clrn(!rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\write2~q ),
	.prn(vcc));
defparam write2.is_wysiwyg = "true";
defparam write2.power_up = "low";

cyclonev_lcell_comb \always2~2 (
	.dataa(!\write1~q ),
	.datab(!\write2~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always2~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always2~2 .extended_lut = "off";
defparam \always2~2 .lut_mask = 64'h6666666666666666;
defparam \always2~2 .shared_arith = "off";

dffeas write_valid(
	.clk(altera_internal_jtag),
	.d(\td_shift[10]~q ),
	.asdata(vcc),
	.clrn(!clr_reg),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_stalled~1_combout ),
	.q(\write_valid~q ),
	.prn(vcc));
defparam write_valid.is_wysiwyg = "true";
defparam write_valid.power_up = "low";

cyclonev_lcell_comb \t_pause~0 (
	.dataa(!t_dav),
	.datab(!\write_stalled~q ),
	.datac(!\rst2~q ),
	.datad(!\always2~1_combout ),
	.datae(!\always2~2_combout ),
	.dataf(!\write_valid~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\t_pause~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \t_pause~0 .extended_lut = "off";
defparam \t_pause~0 .lut_mask = 64'hFFFFFFFF7FFFFFFF;
defparam \t_pause~0 .shared_arith = "off";

cyclonev_lcell_comb \t_ena~0 (
	.dataa(!t_dav),
	.datab(!\write_stalled~q ),
	.datac(!\rst2~q ),
	.datad(!t_ena1),
	.datae(!\always2~2_combout ),
	.dataf(!\write_valid~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\t_ena~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \t_ena~0 .extended_lut = "off";
defparam \t_ena~0 .lut_mask = 64'hEFFFFFFFFFFFFFFF;
defparam \t_ena~0 .shared_arith = "off";

endmodule

module processor_processor_jtag_uart_scfifo_r (
	q_b_0,
	q_b_5,
	q_b_4,
	q_b_6,
	q_b_7,
	q_b_3,
	q_b_2,
	q_b_1,
	r_sync_rst,
	b_full,
	counter_reg_bit_0,
	counter_reg_bit_5,
	counter_reg_bit_4,
	b_non_empty,
	counter_reg_bit_3,
	counter_reg_bit_2,
	counter_reg_bit_1,
	fifo_rd,
	t_ena,
	wr_rfifo,
	wdata_0,
	wdata_5,
	wdata_4,
	wdata_6,
	wdata_7,
	wdata_3,
	wdata_2,
	wdata_1,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_0;
output 	q_b_5;
output 	q_b_4;
output 	q_b_6;
output 	q_b_7;
output 	q_b_3;
output 	q_b_2;
output 	q_b_1;
input 	r_sync_rst;
output 	b_full;
output 	counter_reg_bit_0;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
output 	b_non_empty;
output 	counter_reg_bit_3;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
input 	fifo_rd;
input 	t_ena;
input 	wr_rfifo;
input 	wdata_0;
input 	wdata_5;
input 	wdata_4;
input 	wdata_6;
input 	wdata_7;
input 	wdata_3;
input 	wdata_2;
input 	wdata_1;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



processor_scfifo_1 rfifo(
	.q({q_b_7,q_b_6,q_b_5,q_b_4,q_b_3,q_b_2,q_b_1,q_b_0}),
	.r_sync_rst(r_sync_rst),
	.b_full(b_full),
	.counter_reg_bit_0(counter_reg_bit_0),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_4(counter_reg_bit_4),
	.b_non_empty(b_non_empty),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_1(counter_reg_bit_1),
	.fifo_rd(fifo_rd),
	.t_ena(t_ena),
	.wrreq(wr_rfifo),
	.data({wdata_7,wdata_6,wdata_5,wdata_4,wdata_3,wdata_2,wdata_1,wdata_0}),
	.clock(clk_clk));

endmodule

module processor_scfifo_1 (
	q,
	r_sync_rst,
	b_full,
	counter_reg_bit_0,
	counter_reg_bit_5,
	counter_reg_bit_4,
	b_non_empty,
	counter_reg_bit_3,
	counter_reg_bit_2,
	counter_reg_bit_1,
	fifo_rd,
	t_ena,
	wrreq,
	data,
	clock)/* synthesis synthesis_greybox=1 */;
output 	[7:0] q;
input 	r_sync_rst;
output 	b_full;
output 	counter_reg_bit_0;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
output 	b_non_empty;
output 	counter_reg_bit_3;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
input 	fifo_rd;
input 	t_ena;
input 	wrreq;
input 	[7:0] data;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



processor_scfifo_3291 auto_generated(
	.q({q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.r_sync_rst(r_sync_rst),
	.b_full(b_full),
	.counter_reg_bit_0(counter_reg_bit_0),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_4(counter_reg_bit_4),
	.b_non_empty(b_non_empty),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_1(counter_reg_bit_1),
	.fifo_rd(fifo_rd),
	.t_ena(t_ena),
	.wrreq(wrreq),
	.data({data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.clock(clock));

endmodule

module processor_scfifo_3291 (
	q,
	r_sync_rst,
	b_full,
	counter_reg_bit_0,
	counter_reg_bit_5,
	counter_reg_bit_4,
	b_non_empty,
	counter_reg_bit_3,
	counter_reg_bit_2,
	counter_reg_bit_1,
	fifo_rd,
	t_ena,
	wrreq,
	data,
	clock)/* synthesis synthesis_greybox=1 */;
output 	[7:0] q;
input 	r_sync_rst;
output 	b_full;
output 	counter_reg_bit_0;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
output 	b_non_empty;
output 	counter_reg_bit_3;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
input 	fifo_rd;
input 	t_ena;
input 	wrreq;
input 	[7:0] data;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



processor_a_dpfifo_5771 dpfifo(
	.q({q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.r_sync_rst(r_sync_rst),
	.b_full(b_full),
	.counter_reg_bit_0(counter_reg_bit_0),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_4(counter_reg_bit_4),
	.b_non_empty(b_non_empty),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_1(counter_reg_bit_1),
	.fifo_rd(fifo_rd),
	.t_ena(t_ena),
	.wreq(wrreq),
	.data({data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.clock(clock));

endmodule

module processor_a_dpfifo_5771 (
	q,
	r_sync_rst,
	b_full,
	counter_reg_bit_0,
	counter_reg_bit_5,
	counter_reg_bit_4,
	b_non_empty,
	counter_reg_bit_3,
	counter_reg_bit_2,
	counter_reg_bit_1,
	fifo_rd,
	t_ena,
	wreq,
	data,
	clock)/* synthesis synthesis_greybox=1 */;
output 	[7:0] q;
input 	r_sync_rst;
output 	b_full;
output 	counter_reg_bit_0;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
output 	b_non_empty;
output 	counter_reg_bit_3;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
input 	fifo_rd;
input 	t_ena;
input 	wreq;
input 	[7:0] data;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \wr_ptr|counter_reg_bit[0]~q ;
wire \wr_ptr|counter_reg_bit[1]~q ;
wire \wr_ptr|counter_reg_bit[2]~q ;
wire \wr_ptr|counter_reg_bit[3]~q ;
wire \wr_ptr|counter_reg_bit[4]~q ;
wire \wr_ptr|counter_reg_bit[5]~q ;
wire \rd_ptr_count|counter_reg_bit[0]~q ;
wire \rd_ptr_count|counter_reg_bit[1]~q ;
wire \rd_ptr_count|counter_reg_bit[2]~q ;
wire \rd_ptr_count|counter_reg_bit[3]~q ;
wire \rd_ptr_count|counter_reg_bit[4]~q ;
wire \rd_ptr_count|counter_reg_bit[5]~q ;


processor_a_fefifo_7cf fifo_state(
	.r_sync_rst(r_sync_rst),
	.b_full1(b_full),
	.counter_reg_bit_0(counter_reg_bit_0),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_4(counter_reg_bit_4),
	.b_non_empty1(b_non_empty),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_1(counter_reg_bit_1),
	.fifo_rd(fifo_rd),
	.t_ena(t_ena),
	.wr_rfifo(wreq),
	.clock(clock));

processor_cntr_jgb_1 wr_ptr(
	.r_sync_rst(r_sync_rst),
	.wr_rfifo(wreq),
	.counter_reg_bit_0(\wr_ptr|counter_reg_bit[0]~q ),
	.counter_reg_bit_1(\wr_ptr|counter_reg_bit[1]~q ),
	.counter_reg_bit_2(\wr_ptr|counter_reg_bit[2]~q ),
	.counter_reg_bit_3(\wr_ptr|counter_reg_bit[3]~q ),
	.counter_reg_bit_4(\wr_ptr|counter_reg_bit[4]~q ),
	.counter_reg_bit_5(\wr_ptr|counter_reg_bit[5]~q ),
	.clock(clock));

processor_cntr_jgb rd_ptr_count(
	.r_sync_rst(r_sync_rst),
	.fifo_rd(fifo_rd),
	.counter_reg_bit_0(\rd_ptr_count|counter_reg_bit[0]~q ),
	.counter_reg_bit_1(\rd_ptr_count|counter_reg_bit[1]~q ),
	.counter_reg_bit_2(\rd_ptr_count|counter_reg_bit[2]~q ),
	.counter_reg_bit_3(\rd_ptr_count|counter_reg_bit[3]~q ),
	.counter_reg_bit_4(\rd_ptr_count|counter_reg_bit[4]~q ),
	.counter_reg_bit_5(\rd_ptr_count|counter_reg_bit[5]~q ),
	.clock(clock));

processor_altsyncram_7pu1 FIFOram(
	.q_b({q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.clocken1(fifo_rd),
	.wren_a(wreq),
	.data_a({data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.address_a({\wr_ptr|counter_reg_bit[5]~q ,\wr_ptr|counter_reg_bit[4]~q ,\wr_ptr|counter_reg_bit[3]~q ,\wr_ptr|counter_reg_bit[2]~q ,\wr_ptr|counter_reg_bit[1]~q ,\wr_ptr|counter_reg_bit[0]~q }),
	.address_b({\rd_ptr_count|counter_reg_bit[5]~q ,\rd_ptr_count|counter_reg_bit[4]~q ,\rd_ptr_count|counter_reg_bit[3]~q ,\rd_ptr_count|counter_reg_bit[2]~q ,\rd_ptr_count|counter_reg_bit[1]~q ,\rd_ptr_count|counter_reg_bit[0]~q }),
	.clock1(clock),
	.clock0(clock));

endmodule

module processor_a_fefifo_7cf (
	r_sync_rst,
	b_full1,
	counter_reg_bit_0,
	counter_reg_bit_5,
	counter_reg_bit_4,
	b_non_empty1,
	counter_reg_bit_3,
	counter_reg_bit_2,
	counter_reg_bit_1,
	fifo_rd,
	t_ena,
	wr_rfifo,
	clock)/* synthesis synthesis_greybox=1 */;
input 	r_sync_rst;
output 	b_full1;
output 	counter_reg_bit_0;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
output 	b_non_empty1;
output 	counter_reg_bit_3;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
input 	fifo_rd;
input 	t_ena;
input 	wr_rfifo;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \_~0_combout ;
wire \b_full~0_combout ;
wire \b_full~1_combout ;
wire \_~1_combout ;
wire \_~2_combout ;
wire \b_non_empty~0_combout ;


processor_cntr_vg7 count_usedw(
	.r_sync_rst(r_sync_rst),
	.counter_reg_bit_0(counter_reg_bit_0),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_4(counter_reg_bit_4),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_1(counter_reg_bit_1),
	.wr_rfifo(wr_rfifo),
	._(\_~0_combout ),
	.clock(clock));

cyclonev_lcell_comb \_~0 (
	.dataa(!fifo_rd),
	.datab(!wr_rfifo),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\_~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \_~0 .extended_lut = "off";
defparam \_~0 .lut_mask = 64'h6666666666666666;
defparam \_~0 .shared_arith = "off";

dffeas b_full(
	.clk(clock),
	.d(\b_full~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(b_full1),
	.prn(vcc));
defparam b_full.is_wysiwyg = "true";
defparam b_full.power_up = "low";

dffeas b_non_empty(
	.clk(clock),
	.d(\b_non_empty~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(b_non_empty1),
	.prn(vcc));
defparam b_non_empty.is_wysiwyg = "true";
defparam b_non_empty.power_up = "low";

cyclonev_lcell_comb \b_full~0 (
	.dataa(!counter_reg_bit_3),
	.datab(!counter_reg_bit_2),
	.datac(!counter_reg_bit_5),
	.datad(!counter_reg_bit_4),
	.datae(!b_non_empty1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\b_full~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \b_full~0 .extended_lut = "off";
defparam \b_full~0 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \b_full~0 .shared_arith = "off";

cyclonev_lcell_comb \b_full~1 (
	.dataa(!b_full1),
	.datab(!counter_reg_bit_0),
	.datac(!counter_reg_bit_1),
	.datad(!fifo_rd),
	.datae(!t_ena),
	.dataf(!\b_full~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\b_full~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \b_full~1 .extended_lut = "off";
defparam \b_full~1 .lut_mask = 64'hFF7FFFFFFFFFFFFF;
defparam \b_full~1 .shared_arith = "off";

cyclonev_lcell_comb \_~1 (
	.dataa(!counter_reg_bit_3),
	.datab(!counter_reg_bit_5),
	.datac(!counter_reg_bit_4),
	.datad(!wr_rfifo),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\_~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \_~1 .extended_lut = "off";
defparam \_~1 .lut_mask = 64'hFFFEFFFEFFFEFFFE;
defparam \_~1 .shared_arith = "off";

cyclonev_lcell_comb \_~2 (
	.dataa(!counter_reg_bit_0),
	.datab(!counter_reg_bit_2),
	.datac(!counter_reg_bit_1),
	.datad(!\_~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\_~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \_~2 .extended_lut = "off";
defparam \_~2 .lut_mask = 64'hFDFFFDFFFDFFFDFF;
defparam \_~2 .shared_arith = "off";

cyclonev_lcell_comb \b_non_empty~0 (
	.dataa(!b_full1),
	.datab(!b_non_empty1),
	.datac(!fifo_rd),
	.datad(!t_ena),
	.datae(!\_~2_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\b_non_empty~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \b_non_empty~0 .extended_lut = "off";
defparam \b_non_empty~0 .lut_mask = 64'hF7FFD5FFF7FFD5FF;
defparam \b_non_empty~0 .shared_arith = "off";

endmodule

module processor_cntr_vg7 (
	r_sync_rst,
	counter_reg_bit_0,
	counter_reg_bit_5,
	counter_reg_bit_4,
	counter_reg_bit_3,
	counter_reg_bit_2,
	counter_reg_bit_1,
	wr_rfifo,
	_,
	clock)/* synthesis synthesis_greybox=1 */;
input 	r_sync_rst;
output 	counter_reg_bit_0;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
output 	counter_reg_bit_3;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
input 	wr_rfifo;
input 	_;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~sumout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~COUT ;
wire \counter_comb_bita4~COUT ;
wire \counter_comb_bita5~sumout ;
wire \counter_comb_bita4~sumout ;
wire \counter_comb_bita3~sumout ;
wire \counter_comb_bita2~sumout ;
wire \counter_comb_bita1~sumout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[5] (
	.clk(clock),
	.d(\counter_comb_bita5~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_5),
	.prn(vcc));
defparam \counter_reg_bit[5] .is_wysiwyg = "true";
defparam \counter_reg_bit[5] .power_up = "low";

dffeas \counter_reg_bit[4] (
	.clk(clock),
	.d(\counter_comb_bita4~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_4),
	.prn(vcc));
defparam \counter_reg_bit[4] .is_wysiwyg = "true";
defparam \counter_reg_bit[4] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

cyclonev_lcell_comb counter_comb_bita0(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita0~sumout ),
	.cout(\counter_comb_bita0~COUT ),
	.shareout());
defparam counter_comb_bita0.extended_lut = "off";
defparam counter_comb_bita0.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita0.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita1(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_1),
	.datae(gnd),
	.dataf(!wr_rfifo),
	.datag(gnd),
	.cin(\counter_comb_bita0~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita1~sumout ),
	.cout(\counter_comb_bita1~COUT ),
	.shareout());
defparam counter_comb_bita1.extended_lut = "off";
defparam counter_comb_bita1.lut_mask = 64'h000000FF000000FF;
defparam counter_comb_bita1.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita2(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_2),
	.datae(gnd),
	.dataf(!wr_rfifo),
	.datag(gnd),
	.cin(\counter_comb_bita1~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita2~sumout ),
	.cout(\counter_comb_bita2~COUT ),
	.shareout());
defparam counter_comb_bita2.extended_lut = "off";
defparam counter_comb_bita2.lut_mask = 64'h000000FF000000FF;
defparam counter_comb_bita2.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita3(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_3),
	.datae(gnd),
	.dataf(!wr_rfifo),
	.datag(gnd),
	.cin(\counter_comb_bita2~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita3~sumout ),
	.cout(\counter_comb_bita3~COUT ),
	.shareout());
defparam counter_comb_bita3.extended_lut = "off";
defparam counter_comb_bita3.lut_mask = 64'h000000FF000000FF;
defparam counter_comb_bita3.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita4(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_4),
	.datae(gnd),
	.dataf(!wr_rfifo),
	.datag(gnd),
	.cin(\counter_comb_bita3~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita4~sumout ),
	.cout(\counter_comb_bita4~COUT ),
	.shareout());
defparam counter_comb_bita4.extended_lut = "off";
defparam counter_comb_bita4.lut_mask = 64'h000000FF000000FF;
defparam counter_comb_bita4.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita5(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_5),
	.datae(gnd),
	.dataf(!wr_rfifo),
	.datag(gnd),
	.cin(\counter_comb_bita4~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita5~sumout ),
	.cout(),
	.shareout());
defparam counter_comb_bita5.extended_lut = "off";
defparam counter_comb_bita5.lut_mask = 64'h000000FF000000FF;
defparam counter_comb_bita5.shared_arith = "off";

endmodule

module processor_altsyncram_7pu1 (
	q_b,
	clocken1,
	wren_a,
	data_a,
	address_a,
	address_b,
	clock1,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[7:0] q_b;
input 	clocken1;
input 	wren_a;
input 	[7:0] data_a;
input 	[5:0] address_a;
input 	[5:0] address_b;
input 	clock1;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a0_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a4_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;
wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a1_PORTBDATAOUT_bus;

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_b[3] = ram_block1a3_PORTBDATAOUT_bus[0];

assign q_b[2] = ram_block1a2_PORTBDATAOUT_bus[0];

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

cyclonev_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.clk1_core_clock_enable = "ena1";
defparam ram_block1a0.clk1_input_clock_enable = "ena1";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.logical_ram_name = "processor_jtag_uart:jtag_uart|processor_jtag_uart_scfifo_r:the_processor_jtag_uart_scfifo_r|scfifo:rfifo|scfifo_3291:auto_generated|a_dpfifo_5771:dpfifo|altsyncram_7pu1:FIFOram|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a0.operation_mode = "dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 6;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 63;
defparam ram_block1a0.port_a_logical_ram_depth = 64;
defparam ram_block1a0.port_a_logical_ram_width = 8;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_address_clear = "none";
defparam ram_block1a0.port_b_address_clock = "clock1";
defparam ram_block1a0.port_b_address_width = 6;
defparam ram_block1a0.port_b_data_out_clear = "none";
defparam ram_block1a0.port_b_data_out_clock = "none";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 63;
defparam ram_block1a0.port_b_logical_ram_depth = 64;
defparam ram_block1a0.port_b_logical_ram_width = 8;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock1";
defparam ram_block1a0.ram_block_type = "auto";

cyclonev_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a5.clk0_core_clock_enable = "ena0";
defparam ram_block1a5.clk1_core_clock_enable = "ena1";
defparam ram_block1a5.clk1_input_clock_enable = "ena1";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "processor_jtag_uart:jtag_uart|processor_jtag_uart_scfifo_r:the_processor_jtag_uart_scfifo_r|scfifo:rfifo|scfifo_3291:auto_generated|a_dpfifo_5771:dpfifo|altsyncram_7pu1:FIFOram|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 6;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 63;
defparam ram_block1a5.port_a_logical_ram_depth = 64;
defparam ram_block1a5.port_a_logical_ram_width = 8;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_address_clear = "none";
defparam ram_block1a5.port_b_address_clock = "clock1";
defparam ram_block1a5.port_b_address_width = 6;
defparam ram_block1a5.port_b_data_out_clear = "none";
defparam ram_block1a5.port_b_data_out_clock = "none";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 63;
defparam ram_block1a5.port_b_logical_ram_depth = 64;
defparam ram_block1a5.port_b_logical_ram_width = 8;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock1";
defparam ram_block1a5.ram_block_type = "auto";

cyclonev_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a4.clk0_core_clock_enable = "ena0";
defparam ram_block1a4.clk1_core_clock_enable = "ena1";
defparam ram_block1a4.clk1_input_clock_enable = "ena1";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.logical_ram_name = "processor_jtag_uart:jtag_uart|processor_jtag_uart_scfifo_r:the_processor_jtag_uart_scfifo_r|scfifo:rfifo|scfifo_3291:auto_generated|a_dpfifo_5771:dpfifo|altsyncram_7pu1:FIFOram|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a4.operation_mode = "dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 6;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 63;
defparam ram_block1a4.port_a_logical_ram_depth = 64;
defparam ram_block1a4.port_a_logical_ram_width = 8;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_address_clear = "none";
defparam ram_block1a4.port_b_address_clock = "clock1";
defparam ram_block1a4.port_b_address_width = 6;
defparam ram_block1a4.port_b_data_out_clear = "none";
defparam ram_block1a4.port_b_data_out_clock = "none";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 63;
defparam ram_block1a4.port_b_logical_ram_depth = 64;
defparam ram_block1a4.port_b_logical_ram_width = 8;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock1";
defparam ram_block1a4.ram_block_type = "auto";

cyclonev_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a6.clk0_core_clock_enable = "ena0";
defparam ram_block1a6.clk1_core_clock_enable = "ena1";
defparam ram_block1a6.clk1_input_clock_enable = "ena1";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "processor_jtag_uart:jtag_uart|processor_jtag_uart_scfifo_r:the_processor_jtag_uart_scfifo_r|scfifo:rfifo|scfifo_3291:auto_generated|a_dpfifo_5771:dpfifo|altsyncram_7pu1:FIFOram|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 6;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 63;
defparam ram_block1a6.port_a_logical_ram_depth = 64;
defparam ram_block1a6.port_a_logical_ram_width = 8;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_address_clear = "none";
defparam ram_block1a6.port_b_address_clock = "clock1";
defparam ram_block1a6.port_b_address_width = 6;
defparam ram_block1a6.port_b_data_out_clear = "none";
defparam ram_block1a6.port_b_data_out_clock = "none";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 63;
defparam ram_block1a6.port_b_logical_ram_depth = 64;
defparam ram_block1a6.port_b_logical_ram_width = 8;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock1";
defparam ram_block1a6.ram_block_type = "auto";

cyclonev_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a7.clk0_core_clock_enable = "ena0";
defparam ram_block1a7.clk1_core_clock_enable = "ena1";
defparam ram_block1a7.clk1_input_clock_enable = "ena1";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "processor_jtag_uart:jtag_uart|processor_jtag_uart_scfifo_r:the_processor_jtag_uart_scfifo_r|scfifo:rfifo|scfifo_3291:auto_generated|a_dpfifo_5771:dpfifo|altsyncram_7pu1:FIFOram|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 6;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 63;
defparam ram_block1a7.port_a_logical_ram_depth = 64;
defparam ram_block1a7.port_a_logical_ram_width = 8;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_address_clear = "none";
defparam ram_block1a7.port_b_address_clock = "clock1";
defparam ram_block1a7.port_b_address_width = 6;
defparam ram_block1a7.port_b_data_out_clear = "none";
defparam ram_block1a7.port_b_data_out_clock = "none";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 63;
defparam ram_block1a7.port_b_logical_ram_depth = 64;
defparam ram_block1a7.port_b_logical_ram_width = 8;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock1";
defparam ram_block1a7.ram_block_type = "auto";

cyclonev_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a3.clk0_core_clock_enable = "ena0";
defparam ram_block1a3.clk1_core_clock_enable = "ena1";
defparam ram_block1a3.clk1_input_clock_enable = "ena1";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.logical_ram_name = "processor_jtag_uart:jtag_uart|processor_jtag_uart_scfifo_r:the_processor_jtag_uart_scfifo_r|scfifo:rfifo|scfifo_3291:auto_generated|a_dpfifo_5771:dpfifo|altsyncram_7pu1:FIFOram|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a3.operation_mode = "dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 6;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 63;
defparam ram_block1a3.port_a_logical_ram_depth = 64;
defparam ram_block1a3.port_a_logical_ram_width = 8;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_address_clear = "none";
defparam ram_block1a3.port_b_address_clock = "clock1";
defparam ram_block1a3.port_b_address_width = 6;
defparam ram_block1a3.port_b_data_out_clear = "none";
defparam ram_block1a3.port_b_data_out_clock = "none";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 63;
defparam ram_block1a3.port_b_logical_ram_depth = 64;
defparam ram_block1a3.port_b_logical_ram_width = 8;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock1";
defparam ram_block1a3.ram_block_type = "auto";

cyclonev_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a2.clk0_core_clock_enable = "ena0";
defparam ram_block1a2.clk1_core_clock_enable = "ena1";
defparam ram_block1a2.clk1_input_clock_enable = "ena1";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.logical_ram_name = "processor_jtag_uart:jtag_uart|processor_jtag_uart_scfifo_r:the_processor_jtag_uart_scfifo_r|scfifo:rfifo|scfifo_3291:auto_generated|a_dpfifo_5771:dpfifo|altsyncram_7pu1:FIFOram|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a2.operation_mode = "dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 6;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 63;
defparam ram_block1a2.port_a_logical_ram_depth = 64;
defparam ram_block1a2.port_a_logical_ram_width = 8;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_address_clear = "none";
defparam ram_block1a2.port_b_address_clock = "clock1";
defparam ram_block1a2.port_b_address_width = 6;
defparam ram_block1a2.port_b_data_out_clear = "none";
defparam ram_block1a2.port_b_data_out_clock = "none";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 63;
defparam ram_block1a2.port_b_logical_ram_depth = 64;
defparam ram_block1a2.port_b_logical_ram_width = 8;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock1";
defparam ram_block1a2.ram_block_type = "auto";

cyclonev_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a1.clk0_core_clock_enable = "ena0";
defparam ram_block1a1.clk1_core_clock_enable = "ena1";
defparam ram_block1a1.clk1_input_clock_enable = "ena1";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.logical_ram_name = "processor_jtag_uart:jtag_uart|processor_jtag_uart_scfifo_r:the_processor_jtag_uart_scfifo_r|scfifo:rfifo|scfifo_3291:auto_generated|a_dpfifo_5771:dpfifo|altsyncram_7pu1:FIFOram|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a1.operation_mode = "dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 6;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 63;
defparam ram_block1a1.port_a_logical_ram_depth = 64;
defparam ram_block1a1.port_a_logical_ram_width = 8;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_address_clear = "none";
defparam ram_block1a1.port_b_address_clock = "clock1";
defparam ram_block1a1.port_b_address_width = 6;
defparam ram_block1a1.port_b_data_out_clear = "none";
defparam ram_block1a1.port_b_data_out_clock = "none";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 63;
defparam ram_block1a1.port_b_logical_ram_depth = 64;
defparam ram_block1a1.port_b_logical_ram_width = 8;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock1";
defparam ram_block1a1.ram_block_type = "auto";

endmodule

module processor_cntr_jgb (
	r_sync_rst,
	fifo_rd,
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_2,
	counter_reg_bit_3,
	counter_reg_bit_4,
	counter_reg_bit_5,
	clock)/* synthesis synthesis_greybox=1 */;
input 	r_sync_rst;
input 	fifo_rd;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_2;
output 	counter_reg_bit_3;
output 	counter_reg_bit_4;
output 	counter_reg_bit_5;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~sumout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~sumout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~sumout ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~sumout ;
wire \counter_comb_bita3~COUT ;
wire \counter_comb_bita4~sumout ;
wire \counter_comb_bita4~COUT ;
wire \counter_comb_bita5~sumout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fifo_rd),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fifo_rd),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fifo_rd),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fifo_rd),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

dffeas \counter_reg_bit[4] (
	.clk(clock),
	.d(\counter_comb_bita4~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fifo_rd),
	.q(counter_reg_bit_4),
	.prn(vcc));
defparam \counter_reg_bit[4] .is_wysiwyg = "true";
defparam \counter_reg_bit[4] .power_up = "low";

dffeas \counter_reg_bit[5] (
	.clk(clock),
	.d(\counter_comb_bita5~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fifo_rd),
	.q(counter_reg_bit_5),
	.prn(vcc));
defparam \counter_reg_bit[5] .is_wysiwyg = "true";
defparam \counter_reg_bit[5] .power_up = "low";

cyclonev_lcell_comb counter_comb_bita0(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita0~sumout ),
	.cout(\counter_comb_bita0~COUT ),
	.shareout());
defparam counter_comb_bita0.extended_lut = "off";
defparam counter_comb_bita0.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita0.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita1(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita0~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita1~sumout ),
	.cout(\counter_comb_bita1~COUT ),
	.shareout());
defparam counter_comb_bita1.extended_lut = "off";
defparam counter_comb_bita1.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita1.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita2(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita1~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita2~sumout ),
	.cout(\counter_comb_bita2~COUT ),
	.shareout());
defparam counter_comb_bita2.extended_lut = "off";
defparam counter_comb_bita2.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita2.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita3(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita2~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita3~sumout ),
	.cout(\counter_comb_bita3~COUT ),
	.shareout());
defparam counter_comb_bita3.extended_lut = "off";
defparam counter_comb_bita3.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita3.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita4(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_4),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita3~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita4~sumout ),
	.cout(\counter_comb_bita4~COUT ),
	.shareout());
defparam counter_comb_bita4.extended_lut = "off";
defparam counter_comb_bita4.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita4.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita5(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_5),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita4~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita5~sumout ),
	.cout(),
	.shareout());
defparam counter_comb_bita5.extended_lut = "off";
defparam counter_comb_bita5.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita5.shared_arith = "off";

endmodule

module processor_cntr_jgb_1 (
	r_sync_rst,
	wr_rfifo,
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_2,
	counter_reg_bit_3,
	counter_reg_bit_4,
	counter_reg_bit_5,
	clock)/* synthesis synthesis_greybox=1 */;
input 	r_sync_rst;
input 	wr_rfifo;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_2;
output 	counter_reg_bit_3;
output 	counter_reg_bit_4;
output 	counter_reg_bit_5;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~sumout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~sumout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~sumout ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~sumout ;
wire \counter_comb_bita3~COUT ;
wire \counter_comb_bita4~sumout ;
wire \counter_comb_bita4~COUT ;
wire \counter_comb_bita5~sumout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wr_rfifo),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wr_rfifo),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wr_rfifo),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wr_rfifo),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

dffeas \counter_reg_bit[4] (
	.clk(clock),
	.d(\counter_comb_bita4~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wr_rfifo),
	.q(counter_reg_bit_4),
	.prn(vcc));
defparam \counter_reg_bit[4] .is_wysiwyg = "true";
defparam \counter_reg_bit[4] .power_up = "low";

dffeas \counter_reg_bit[5] (
	.clk(clock),
	.d(\counter_comb_bita5~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(wr_rfifo),
	.q(counter_reg_bit_5),
	.prn(vcc));
defparam \counter_reg_bit[5] .is_wysiwyg = "true";
defparam \counter_reg_bit[5] .power_up = "low";

cyclonev_lcell_comb counter_comb_bita0(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita0~sumout ),
	.cout(\counter_comb_bita0~COUT ),
	.shareout());
defparam counter_comb_bita0.extended_lut = "off";
defparam counter_comb_bita0.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita0.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita1(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita0~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita1~sumout ),
	.cout(\counter_comb_bita1~COUT ),
	.shareout());
defparam counter_comb_bita1.extended_lut = "off";
defparam counter_comb_bita1.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita1.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita2(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita1~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita2~sumout ),
	.cout(\counter_comb_bita2~COUT ),
	.shareout());
defparam counter_comb_bita2.extended_lut = "off";
defparam counter_comb_bita2.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita2.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita3(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita2~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita3~sumout ),
	.cout(\counter_comb_bita3~COUT ),
	.shareout());
defparam counter_comb_bita3.extended_lut = "off";
defparam counter_comb_bita3.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita3.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita4(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_4),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita3~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita4~sumout ),
	.cout(\counter_comb_bita4~COUT ),
	.shareout());
defparam counter_comb_bita4.extended_lut = "off";
defparam counter_comb_bita4.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita4.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita5(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_5),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita4~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita5~sumout ),
	.cout(),
	.shareout());
defparam counter_comb_bita5.extended_lut = "off";
defparam counter_comb_bita5.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita5.shared_arith = "off";

endmodule

module processor_processor_jtag_uart_scfifo_w (
	q_b_7,
	q_b_0,
	q_b_1,
	q_b_2,
	q_b_3,
	q_b_6,
	q_b_5,
	q_b_4,
	M_st_data_0,
	r_sync_rst,
	M_st_data_1,
	M_st_data_2,
	M_st_data_3,
	M_st_data_4,
	M_st_data_5,
	M_st_data_6,
	M_st_data_7,
	b_full,
	counter_reg_bit_5,
	counter_reg_bit_4,
	counter_reg_bit_0,
	counter_reg_bit_3,
	counter_reg_bit_2,
	counter_reg_bit_1,
	fifo_wr,
	b_non_empty,
	r_val,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_7;
output 	q_b_0;
output 	q_b_1;
output 	q_b_2;
output 	q_b_3;
output 	q_b_6;
output 	q_b_5;
output 	q_b_4;
input 	M_st_data_0;
input 	r_sync_rst;
input 	M_st_data_1;
input 	M_st_data_2;
input 	M_st_data_3;
input 	M_st_data_4;
input 	M_st_data_5;
input 	M_st_data_6;
input 	M_st_data_7;
output 	b_full;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
output 	counter_reg_bit_0;
output 	counter_reg_bit_3;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
input 	fifo_wr;
output 	b_non_empty;
input 	r_val;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



processor_scfifo_2 wfifo(
	.q({q_b_7,q_b_6,q_b_5,q_b_4,q_b_3,q_b_2,q_b_1,q_b_0}),
	.data({M_st_data_7,M_st_data_6,M_st_data_5,M_st_data_4,M_st_data_3,M_st_data_2,M_st_data_1,M_st_data_0}),
	.r_sync_rst(r_sync_rst),
	.b_full(b_full),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_4(counter_reg_bit_4),
	.counter_reg_bit_0(counter_reg_bit_0),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_1(counter_reg_bit_1),
	.wrreq(fifo_wr),
	.b_non_empty(b_non_empty),
	.r_val(r_val),
	.clock(clk_clk));

endmodule

module processor_scfifo_2 (
	q,
	data,
	r_sync_rst,
	b_full,
	counter_reg_bit_5,
	counter_reg_bit_4,
	counter_reg_bit_0,
	counter_reg_bit_3,
	counter_reg_bit_2,
	counter_reg_bit_1,
	wrreq,
	b_non_empty,
	r_val,
	clock)/* synthesis synthesis_greybox=1 */;
output 	[7:0] q;
input 	[7:0] data;
input 	r_sync_rst;
output 	b_full;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
output 	counter_reg_bit_0;
output 	counter_reg_bit_3;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
input 	wrreq;
output 	b_non_empty;
input 	r_val;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



processor_scfifo_3291_1 auto_generated(
	.q({q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.data({data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.r_sync_rst(r_sync_rst),
	.b_full(b_full),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_4(counter_reg_bit_4),
	.counter_reg_bit_0(counter_reg_bit_0),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_1(counter_reg_bit_1),
	.wrreq(wrreq),
	.b_non_empty(b_non_empty),
	.r_val(r_val),
	.clock(clock));

endmodule

module processor_scfifo_3291_1 (
	q,
	data,
	r_sync_rst,
	b_full,
	counter_reg_bit_5,
	counter_reg_bit_4,
	counter_reg_bit_0,
	counter_reg_bit_3,
	counter_reg_bit_2,
	counter_reg_bit_1,
	wrreq,
	b_non_empty,
	r_val,
	clock)/* synthesis synthesis_greybox=1 */;
output 	[7:0] q;
input 	[7:0] data;
input 	r_sync_rst;
output 	b_full;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
output 	counter_reg_bit_0;
output 	counter_reg_bit_3;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
input 	wrreq;
output 	b_non_empty;
input 	r_val;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



processor_a_dpfifo_5771_1 dpfifo(
	.q({q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.data({data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.r_sync_rst(r_sync_rst),
	.b_full(b_full),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_4(counter_reg_bit_4),
	.counter_reg_bit_0(counter_reg_bit_0),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_1(counter_reg_bit_1),
	.wreq(wrreq),
	.b_non_empty(b_non_empty),
	.r_val(r_val),
	.clock(clock));

endmodule

module processor_a_dpfifo_5771_1 (
	q,
	data,
	r_sync_rst,
	b_full,
	counter_reg_bit_5,
	counter_reg_bit_4,
	counter_reg_bit_0,
	counter_reg_bit_3,
	counter_reg_bit_2,
	counter_reg_bit_1,
	wreq,
	b_non_empty,
	r_val,
	clock)/* synthesis synthesis_greybox=1 */;
output 	[7:0] q;
input 	[7:0] data;
input 	r_sync_rst;
output 	b_full;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
output 	counter_reg_bit_0;
output 	counter_reg_bit_3;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
input 	wreq;
output 	b_non_empty;
input 	r_val;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \wr_ptr|counter_reg_bit[0]~q ;
wire \wr_ptr|counter_reg_bit[1]~q ;
wire \wr_ptr|counter_reg_bit[2]~q ;
wire \wr_ptr|counter_reg_bit[3]~q ;
wire \wr_ptr|counter_reg_bit[4]~q ;
wire \wr_ptr|counter_reg_bit[5]~q ;
wire \rd_ptr_count|counter_reg_bit[0]~q ;
wire \rd_ptr_count|counter_reg_bit[1]~q ;
wire \rd_ptr_count|counter_reg_bit[2]~q ;
wire \rd_ptr_count|counter_reg_bit[3]~q ;
wire \rd_ptr_count|counter_reg_bit[4]~q ;
wire \rd_ptr_count|counter_reg_bit[5]~q ;


processor_cntr_jgb_3 wr_ptr(
	.r_sync_rst(r_sync_rst),
	.fifo_wr(wreq),
	.counter_reg_bit_0(\wr_ptr|counter_reg_bit[0]~q ),
	.counter_reg_bit_1(\wr_ptr|counter_reg_bit[1]~q ),
	.counter_reg_bit_2(\wr_ptr|counter_reg_bit[2]~q ),
	.counter_reg_bit_3(\wr_ptr|counter_reg_bit[3]~q ),
	.counter_reg_bit_4(\wr_ptr|counter_reg_bit[4]~q ),
	.counter_reg_bit_5(\wr_ptr|counter_reg_bit[5]~q ),
	.clock(clock));

processor_cntr_jgb_2 rd_ptr_count(
	.r_sync_rst(r_sync_rst),
	.r_val(r_val),
	.counter_reg_bit_0(\rd_ptr_count|counter_reg_bit[0]~q ),
	.counter_reg_bit_1(\rd_ptr_count|counter_reg_bit[1]~q ),
	.counter_reg_bit_2(\rd_ptr_count|counter_reg_bit[2]~q ),
	.counter_reg_bit_3(\rd_ptr_count|counter_reg_bit[3]~q ),
	.counter_reg_bit_4(\rd_ptr_count|counter_reg_bit[4]~q ),
	.counter_reg_bit_5(\rd_ptr_count|counter_reg_bit[5]~q ),
	.clock(clock));

processor_altsyncram_7pu1_1 FIFOram(
	.q_b({q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0]}),
	.data_a({data[7],data[6],data[5],data[4],data[3],data[2],data[1],data[0]}),
	.wren_a(wreq),
	.clocken1(r_val),
	.address_a({\wr_ptr|counter_reg_bit[5]~q ,\wr_ptr|counter_reg_bit[4]~q ,\wr_ptr|counter_reg_bit[3]~q ,\wr_ptr|counter_reg_bit[2]~q ,\wr_ptr|counter_reg_bit[1]~q ,\wr_ptr|counter_reg_bit[0]~q }),
	.address_b({\rd_ptr_count|counter_reg_bit[5]~q ,\rd_ptr_count|counter_reg_bit[4]~q ,\rd_ptr_count|counter_reg_bit[3]~q ,\rd_ptr_count|counter_reg_bit[2]~q ,\rd_ptr_count|counter_reg_bit[1]~q ,\rd_ptr_count|counter_reg_bit[0]~q }),
	.clock1(clock),
	.clock0(clock));

processor_a_fefifo_7cf_1 fifo_state(
	.r_sync_rst(r_sync_rst),
	.b_full1(b_full),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_4(counter_reg_bit_4),
	.counter_reg_bit_0(counter_reg_bit_0),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_1(counter_reg_bit_1),
	.fifo_wr(wreq),
	.b_non_empty1(b_non_empty),
	.r_val(r_val),
	.clock(clock));

endmodule

module processor_a_fefifo_7cf_1 (
	r_sync_rst,
	b_full1,
	counter_reg_bit_5,
	counter_reg_bit_4,
	counter_reg_bit_0,
	counter_reg_bit_3,
	counter_reg_bit_2,
	counter_reg_bit_1,
	fifo_wr,
	b_non_empty1,
	r_val,
	clock)/* synthesis synthesis_greybox=1 */;
input 	r_sync_rst;
output 	b_full1;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
output 	counter_reg_bit_0;
output 	counter_reg_bit_3;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
input 	fifo_wr;
output 	b_non_empty1;
input 	r_val;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \_~0_combout ;
wire \b_full~0_combout ;
wire \b_full~1_combout ;
wire \b_non_empty~0_combout ;
wire \b_non_empty~1_combout ;
wire \b_non_empty~2_combout ;


processor_cntr_vg7_1 count_usedw(
	.r_sync_rst(r_sync_rst),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_4(counter_reg_bit_4),
	.counter_reg_bit_0(counter_reg_bit_0),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_1(counter_reg_bit_1),
	.fifo_wr(fifo_wr),
	._(\_~0_combout ),
	.clock(clock));

cyclonev_lcell_comb \_~0 (
	.dataa(!fifo_wr),
	.datab(!r_val),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\_~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \_~0 .extended_lut = "off";
defparam \_~0 .lut_mask = 64'h6666666666666666;
defparam \_~0 .shared_arith = "off";

dffeas b_full(
	.clk(clock),
	.d(\b_full~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(b_full1),
	.prn(vcc));
defparam b_full.is_wysiwyg = "true";
defparam b_full.power_up = "low";

dffeas b_non_empty(
	.clk(clock),
	.d(\b_non_empty~2_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(b_non_empty1),
	.prn(vcc));
defparam b_non_empty.is_wysiwyg = "true";
defparam b_non_empty.power_up = "low";

cyclonev_lcell_comb \b_full~0 (
	.dataa(!counter_reg_bit_3),
	.datab(!counter_reg_bit_5),
	.datac(!counter_reg_bit_4),
	.datad(!fifo_wr),
	.datae(!b_non_empty1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\b_full~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \b_full~0 .extended_lut = "off";
defparam \b_full~0 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \b_full~0 .shared_arith = "off";

cyclonev_lcell_comb \b_full~1 (
	.dataa(!counter_reg_bit_0),
	.datab(!counter_reg_bit_2),
	.datac(!counter_reg_bit_1),
	.datad(!b_full1),
	.datae(!r_val),
	.dataf(!\b_full~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\b_full~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \b_full~1 .extended_lut = "off";
defparam \b_full~1 .lut_mask = 64'hFFFF7FFFFFFFFFFF;
defparam \b_full~1 .shared_arith = "off";

cyclonev_lcell_comb \b_non_empty~0 (
	.dataa(!counter_reg_bit_2),
	.datab(!counter_reg_bit_1),
	.datac(!counter_reg_bit_5),
	.datad(!counter_reg_bit_4),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\b_non_empty~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \b_non_empty~0 .extended_lut = "off";
defparam \b_non_empty~0 .lut_mask = 64'hFFFEFFFEFFFEFFFE;
defparam \b_non_empty~0 .shared_arith = "off";

cyclonev_lcell_comb \b_non_empty~1 (
	.dataa(!counter_reg_bit_0),
	.datab(!counter_reg_bit_3),
	.datac(!r_val),
	.datad(!\b_non_empty~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\b_non_empty~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \b_non_empty~1 .extended_lut = "off";
defparam \b_non_empty~1 .lut_mask = 64'hDFFFDFFFDFFFDFFF;
defparam \b_non_empty~1 .shared_arith = "off";

cyclonev_lcell_comb \b_non_empty~2 (
	.dataa(!b_full1),
	.datab(!fifo_wr),
	.datac(!b_non_empty1),
	.datad(!\b_non_empty~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\b_non_empty~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \b_non_empty~2 .extended_lut = "off";
defparam \b_non_empty~2 .lut_mask = 64'hFF7FFF7FFF7FFF7F;
defparam \b_non_empty~2 .shared_arith = "off";

endmodule

module processor_cntr_vg7_1 (
	r_sync_rst,
	counter_reg_bit_5,
	counter_reg_bit_4,
	counter_reg_bit_0,
	counter_reg_bit_3,
	counter_reg_bit_2,
	counter_reg_bit_1,
	fifo_wr,
	_,
	clock)/* synthesis synthesis_greybox=1 */;
input 	r_sync_rst;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
output 	counter_reg_bit_0;
output 	counter_reg_bit_3;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
input 	fifo_wr;
input 	_;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~COUT ;
wire \counter_comb_bita4~COUT ;
wire \counter_comb_bita5~sumout ;
wire \counter_comb_bita4~sumout ;
wire \counter_comb_bita0~sumout ;
wire \counter_comb_bita3~sumout ;
wire \counter_comb_bita2~sumout ;
wire \counter_comb_bita1~sumout ;


dffeas \counter_reg_bit[5] (
	.clk(clock),
	.d(\counter_comb_bita5~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_5),
	.prn(vcc));
defparam \counter_reg_bit[5] .is_wysiwyg = "true";
defparam \counter_reg_bit[5] .power_up = "low";

dffeas \counter_reg_bit[4] (
	.clk(clock),
	.d(\counter_comb_bita4~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_4),
	.prn(vcc));
defparam \counter_reg_bit[4] .is_wysiwyg = "true";
defparam \counter_reg_bit[4] .power_up = "low";

dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(_),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

cyclonev_lcell_comb counter_comb_bita0(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita0~sumout ),
	.cout(\counter_comb_bita0~COUT ),
	.shareout());
defparam counter_comb_bita0.extended_lut = "off";
defparam counter_comb_bita0.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita0.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita1(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_1),
	.datae(gnd),
	.dataf(!fifo_wr),
	.datag(gnd),
	.cin(\counter_comb_bita0~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita1~sumout ),
	.cout(\counter_comb_bita1~COUT ),
	.shareout());
defparam counter_comb_bita1.extended_lut = "off";
defparam counter_comb_bita1.lut_mask = 64'h000000FF000000FF;
defparam counter_comb_bita1.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita2(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_2),
	.datae(gnd),
	.dataf(!fifo_wr),
	.datag(gnd),
	.cin(\counter_comb_bita1~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita2~sumout ),
	.cout(\counter_comb_bita2~COUT ),
	.shareout());
defparam counter_comb_bita2.extended_lut = "off";
defparam counter_comb_bita2.lut_mask = 64'h000000FF000000FF;
defparam counter_comb_bita2.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita3(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_3),
	.datae(gnd),
	.dataf(!fifo_wr),
	.datag(gnd),
	.cin(\counter_comb_bita2~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita3~sumout ),
	.cout(\counter_comb_bita3~COUT ),
	.shareout());
defparam counter_comb_bita3.extended_lut = "off";
defparam counter_comb_bita3.lut_mask = 64'h000000FF000000FF;
defparam counter_comb_bita3.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita4(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_4),
	.datae(gnd),
	.dataf(!fifo_wr),
	.datag(gnd),
	.cin(\counter_comb_bita3~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita4~sumout ),
	.cout(\counter_comb_bita4~COUT ),
	.shareout());
defparam counter_comb_bita4.extended_lut = "off";
defparam counter_comb_bita4.lut_mask = 64'h000000FF000000FF;
defparam counter_comb_bita4.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita5(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_5),
	.datae(gnd),
	.dataf(!fifo_wr),
	.datag(gnd),
	.cin(\counter_comb_bita4~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita5~sumout ),
	.cout(),
	.shareout());
defparam counter_comb_bita5.extended_lut = "off";
defparam counter_comb_bita5.lut_mask = 64'h000000FF000000FF;
defparam counter_comb_bita5.shared_arith = "off";

endmodule

module processor_altsyncram_7pu1_1 (
	q_b,
	data_a,
	wren_a,
	clocken1,
	address_a,
	address_b,
	clock1,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[7:0] q_b;
input 	[7:0] data_a;
input 	wren_a;
input 	clocken1;
input 	[5:0] address_a;
input 	[5:0] address_b;
input 	clock1;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a0_PORTBDATAOUT_bus;
wire [143:0] ram_block1a1_PORTBDATAOUT_bus;
wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a4_PORTBDATAOUT_bus;

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

assign q_b[2] = ram_block1a2_PORTBDATAOUT_bus[0];

assign q_b[3] = ram_block1a3_PORTBDATAOUT_bus[0];

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];

cyclonev_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a7.clk0_core_clock_enable = "ena0";
defparam ram_block1a7.clk1_core_clock_enable = "ena1";
defparam ram_block1a7.clk1_input_clock_enable = "ena1";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "processor_jtag_uart:jtag_uart|processor_jtag_uart_scfifo_w:the_processor_jtag_uart_scfifo_w|scfifo:wfifo|scfifo_3291:auto_generated|a_dpfifo_5771:dpfifo|altsyncram_7pu1:FIFOram|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 6;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 63;
defparam ram_block1a7.port_a_logical_ram_depth = 64;
defparam ram_block1a7.port_a_logical_ram_width = 8;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_address_clear = "none";
defparam ram_block1a7.port_b_address_clock = "clock1";
defparam ram_block1a7.port_b_address_width = 6;
defparam ram_block1a7.port_b_data_out_clear = "none";
defparam ram_block1a7.port_b_data_out_clock = "none";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 63;
defparam ram_block1a7.port_b_logical_ram_depth = 64;
defparam ram_block1a7.port_b_logical_ram_width = 8;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock1";
defparam ram_block1a7.ram_block_type = "auto";

cyclonev_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.clk1_core_clock_enable = "ena1";
defparam ram_block1a0.clk1_input_clock_enable = "ena1";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.logical_ram_name = "processor_jtag_uart:jtag_uart|processor_jtag_uart_scfifo_w:the_processor_jtag_uart_scfifo_w|scfifo:wfifo|scfifo_3291:auto_generated|a_dpfifo_5771:dpfifo|altsyncram_7pu1:FIFOram|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a0.operation_mode = "dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 6;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 63;
defparam ram_block1a0.port_a_logical_ram_depth = 64;
defparam ram_block1a0.port_a_logical_ram_width = 8;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_address_clear = "none";
defparam ram_block1a0.port_b_address_clock = "clock1";
defparam ram_block1a0.port_b_address_width = 6;
defparam ram_block1a0.port_b_data_out_clear = "none";
defparam ram_block1a0.port_b_data_out_clock = "none";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 63;
defparam ram_block1a0.port_b_logical_ram_depth = 64;
defparam ram_block1a0.port_b_logical_ram_width = 8;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock1";
defparam ram_block1a0.ram_block_type = "auto";

cyclonev_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a1.clk0_core_clock_enable = "ena0";
defparam ram_block1a1.clk1_core_clock_enable = "ena1";
defparam ram_block1a1.clk1_input_clock_enable = "ena1";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.logical_ram_name = "processor_jtag_uart:jtag_uart|processor_jtag_uart_scfifo_w:the_processor_jtag_uart_scfifo_w|scfifo:wfifo|scfifo_3291:auto_generated|a_dpfifo_5771:dpfifo|altsyncram_7pu1:FIFOram|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a1.operation_mode = "dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 6;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 63;
defparam ram_block1a1.port_a_logical_ram_depth = 64;
defparam ram_block1a1.port_a_logical_ram_width = 8;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_address_clear = "none";
defparam ram_block1a1.port_b_address_clock = "clock1";
defparam ram_block1a1.port_b_address_width = 6;
defparam ram_block1a1.port_b_data_out_clear = "none";
defparam ram_block1a1.port_b_data_out_clock = "none";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 63;
defparam ram_block1a1.port_b_logical_ram_depth = 64;
defparam ram_block1a1.port_b_logical_ram_width = 8;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock1";
defparam ram_block1a1.ram_block_type = "auto";

cyclonev_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a2.clk0_core_clock_enable = "ena0";
defparam ram_block1a2.clk1_core_clock_enable = "ena1";
defparam ram_block1a2.clk1_input_clock_enable = "ena1";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.logical_ram_name = "processor_jtag_uart:jtag_uart|processor_jtag_uart_scfifo_w:the_processor_jtag_uart_scfifo_w|scfifo:wfifo|scfifo_3291:auto_generated|a_dpfifo_5771:dpfifo|altsyncram_7pu1:FIFOram|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a2.operation_mode = "dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 6;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 63;
defparam ram_block1a2.port_a_logical_ram_depth = 64;
defparam ram_block1a2.port_a_logical_ram_width = 8;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_address_clear = "none";
defparam ram_block1a2.port_b_address_clock = "clock1";
defparam ram_block1a2.port_b_address_width = 6;
defparam ram_block1a2.port_b_data_out_clear = "none";
defparam ram_block1a2.port_b_data_out_clock = "none";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 63;
defparam ram_block1a2.port_b_logical_ram_depth = 64;
defparam ram_block1a2.port_b_logical_ram_width = 8;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock1";
defparam ram_block1a2.ram_block_type = "auto";

cyclonev_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a3.clk0_core_clock_enable = "ena0";
defparam ram_block1a3.clk1_core_clock_enable = "ena1";
defparam ram_block1a3.clk1_input_clock_enable = "ena1";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.logical_ram_name = "processor_jtag_uart:jtag_uart|processor_jtag_uart_scfifo_w:the_processor_jtag_uart_scfifo_w|scfifo:wfifo|scfifo_3291:auto_generated|a_dpfifo_5771:dpfifo|altsyncram_7pu1:FIFOram|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a3.operation_mode = "dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 6;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 63;
defparam ram_block1a3.port_a_logical_ram_depth = 64;
defparam ram_block1a3.port_a_logical_ram_width = 8;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_address_clear = "none";
defparam ram_block1a3.port_b_address_clock = "clock1";
defparam ram_block1a3.port_b_address_width = 6;
defparam ram_block1a3.port_b_data_out_clear = "none";
defparam ram_block1a3.port_b_data_out_clock = "none";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 63;
defparam ram_block1a3.port_b_logical_ram_depth = 64;
defparam ram_block1a3.port_b_logical_ram_width = 8;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock1";
defparam ram_block1a3.ram_block_type = "auto";

cyclonev_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a6.clk0_core_clock_enable = "ena0";
defparam ram_block1a6.clk1_core_clock_enable = "ena1";
defparam ram_block1a6.clk1_input_clock_enable = "ena1";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "processor_jtag_uart:jtag_uart|processor_jtag_uart_scfifo_w:the_processor_jtag_uart_scfifo_w|scfifo:wfifo|scfifo_3291:auto_generated|a_dpfifo_5771:dpfifo|altsyncram_7pu1:FIFOram|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 6;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 63;
defparam ram_block1a6.port_a_logical_ram_depth = 64;
defparam ram_block1a6.port_a_logical_ram_width = 8;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_address_clear = "none";
defparam ram_block1a6.port_b_address_clock = "clock1";
defparam ram_block1a6.port_b_address_width = 6;
defparam ram_block1a6.port_b_data_out_clear = "none";
defparam ram_block1a6.port_b_data_out_clock = "none";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 63;
defparam ram_block1a6.port_b_logical_ram_depth = 64;
defparam ram_block1a6.port_b_logical_ram_width = 8;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock1";
defparam ram_block1a6.ram_block_type = "auto";

cyclonev_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a5.clk0_core_clock_enable = "ena0";
defparam ram_block1a5.clk1_core_clock_enable = "ena1";
defparam ram_block1a5.clk1_input_clock_enable = "ena1";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "processor_jtag_uart:jtag_uart|processor_jtag_uart_scfifo_w:the_processor_jtag_uart_scfifo_w|scfifo:wfifo|scfifo_3291:auto_generated|a_dpfifo_5771:dpfifo|altsyncram_7pu1:FIFOram|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 6;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 63;
defparam ram_block1a5.port_a_logical_ram_depth = 64;
defparam ram_block1a5.port_a_logical_ram_width = 8;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_address_clear = "none";
defparam ram_block1a5.port_b_address_clock = "clock1";
defparam ram_block1a5.port_b_address_width = 6;
defparam ram_block1a5.port_b_data_out_clear = "none";
defparam ram_block1a5.port_b_data_out_clock = "none";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 63;
defparam ram_block1a5.port_b_logical_ram_depth = 64;
defparam ram_block1a5.port_b_logical_ram_width = 8;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock1";
defparam ram_block1a5.ram_block_type = "auto";

cyclonev_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(wren_a),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a4.clk0_core_clock_enable = "ena0";
defparam ram_block1a4.clk1_core_clock_enable = "ena1";
defparam ram_block1a4.clk1_input_clock_enable = "ena1";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.logical_ram_name = "processor_jtag_uart:jtag_uart|processor_jtag_uart_scfifo_w:the_processor_jtag_uart_scfifo_w|scfifo:wfifo|scfifo_3291:auto_generated|a_dpfifo_5771:dpfifo|altsyncram_7pu1:FIFOram|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a4.operation_mode = "dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 6;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 63;
defparam ram_block1a4.port_a_logical_ram_depth = 64;
defparam ram_block1a4.port_a_logical_ram_width = 8;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_address_clear = "none";
defparam ram_block1a4.port_b_address_clock = "clock1";
defparam ram_block1a4.port_b_address_width = 6;
defparam ram_block1a4.port_b_data_out_clear = "none";
defparam ram_block1a4.port_b_data_out_clock = "none";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 63;
defparam ram_block1a4.port_b_logical_ram_depth = 64;
defparam ram_block1a4.port_b_logical_ram_width = 8;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock1";
defparam ram_block1a4.ram_block_type = "auto";

endmodule

module processor_cntr_jgb_2 (
	r_sync_rst,
	r_val,
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_2,
	counter_reg_bit_3,
	counter_reg_bit_4,
	counter_reg_bit_5,
	clock)/* synthesis synthesis_greybox=1 */;
input 	r_sync_rst;
input 	r_val;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_2;
output 	counter_reg_bit_3;
output 	counter_reg_bit_4;
output 	counter_reg_bit_5;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~sumout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~sumout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~sumout ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~sumout ;
wire \counter_comb_bita3~COUT ;
wire \counter_comb_bita4~sumout ;
wire \counter_comb_bita4~COUT ;
wire \counter_comb_bita5~sumout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(r_val),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(r_val),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(r_val),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(r_val),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

dffeas \counter_reg_bit[4] (
	.clk(clock),
	.d(\counter_comb_bita4~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(r_val),
	.q(counter_reg_bit_4),
	.prn(vcc));
defparam \counter_reg_bit[4] .is_wysiwyg = "true";
defparam \counter_reg_bit[4] .power_up = "low";

dffeas \counter_reg_bit[5] (
	.clk(clock),
	.d(\counter_comb_bita5~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(r_val),
	.q(counter_reg_bit_5),
	.prn(vcc));
defparam \counter_reg_bit[5] .is_wysiwyg = "true";
defparam \counter_reg_bit[5] .power_up = "low";

cyclonev_lcell_comb counter_comb_bita0(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita0~sumout ),
	.cout(\counter_comb_bita0~COUT ),
	.shareout());
defparam counter_comb_bita0.extended_lut = "off";
defparam counter_comb_bita0.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita0.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita1(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita0~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita1~sumout ),
	.cout(\counter_comb_bita1~COUT ),
	.shareout());
defparam counter_comb_bita1.extended_lut = "off";
defparam counter_comb_bita1.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita1.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita2(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita1~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita2~sumout ),
	.cout(\counter_comb_bita2~COUT ),
	.shareout());
defparam counter_comb_bita2.extended_lut = "off";
defparam counter_comb_bita2.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita2.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita3(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita2~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita3~sumout ),
	.cout(\counter_comb_bita3~COUT ),
	.shareout());
defparam counter_comb_bita3.extended_lut = "off";
defparam counter_comb_bita3.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita3.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita4(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_4),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita3~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita4~sumout ),
	.cout(\counter_comb_bita4~COUT ),
	.shareout());
defparam counter_comb_bita4.extended_lut = "off";
defparam counter_comb_bita4.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita4.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita5(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_5),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita4~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita5~sumout ),
	.cout(),
	.shareout());
defparam counter_comb_bita5.extended_lut = "off";
defparam counter_comb_bita5.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita5.shared_arith = "off";

endmodule

module processor_cntr_jgb_3 (
	r_sync_rst,
	fifo_wr,
	counter_reg_bit_0,
	counter_reg_bit_1,
	counter_reg_bit_2,
	counter_reg_bit_3,
	counter_reg_bit_4,
	counter_reg_bit_5,
	clock)/* synthesis synthesis_greybox=1 */;
input 	r_sync_rst;
input 	fifo_wr;
output 	counter_reg_bit_0;
output 	counter_reg_bit_1;
output 	counter_reg_bit_2;
output 	counter_reg_bit_3;
output 	counter_reg_bit_4;
output 	counter_reg_bit_5;
input 	clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~sumout ;
wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~sumout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~sumout ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~sumout ;
wire \counter_comb_bita3~COUT ;
wire \counter_comb_bita4~sumout ;
wire \counter_comb_bita4~COUT ;
wire \counter_comb_bita5~sumout ;


dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fifo_wr),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fifo_wr),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fifo_wr),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fifo_wr),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

dffeas \counter_reg_bit[4] (
	.clk(clock),
	.d(\counter_comb_bita4~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fifo_wr),
	.q(counter_reg_bit_4),
	.prn(vcc));
defparam \counter_reg_bit[4] .is_wysiwyg = "true";
defparam \counter_reg_bit[4] .power_up = "low";

dffeas \counter_reg_bit[5] (
	.clk(clock),
	.d(\counter_comb_bita5~sumout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(fifo_wr),
	.q(counter_reg_bit_5),
	.prn(vcc));
defparam \counter_reg_bit[5] .is_wysiwyg = "true";
defparam \counter_reg_bit[5] .power_up = "low";

cyclonev_lcell_comb counter_comb_bita0(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita0~sumout ),
	.cout(\counter_comb_bita0~COUT ),
	.shareout());
defparam counter_comb_bita0.extended_lut = "off";
defparam counter_comb_bita0.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita0.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita1(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita0~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita1~sumout ),
	.cout(\counter_comb_bita1~COUT ),
	.shareout());
defparam counter_comb_bita1.extended_lut = "off";
defparam counter_comb_bita1.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita1.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita2(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita1~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita2~sumout ),
	.cout(\counter_comb_bita2~COUT ),
	.shareout());
defparam counter_comb_bita2.extended_lut = "off";
defparam counter_comb_bita2.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita2.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita3(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita2~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita3~sumout ),
	.cout(\counter_comb_bita3~COUT ),
	.shareout());
defparam counter_comb_bita3.extended_lut = "off";
defparam counter_comb_bita3.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita3.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita4(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_4),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita3~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita4~sumout ),
	.cout(\counter_comb_bita4~COUT ),
	.shareout());
defparam counter_comb_bita4.extended_lut = "off";
defparam counter_comb_bita4.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita4.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita5(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_5),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita4~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita5~sumout ),
	.cout(),
	.shareout());
defparam counter_comb_bita5.extended_lut = "off";
defparam counter_comb_bita5.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita5.shared_arith = "off";

endmodule

module processor_processor_led_pio (
	writedata,
	data_out_0,
	data_out_1,
	data_out_2,
	data_out_3,
	data_out_4,
	data_out_5,
	data_out_6,
	data_out_7,
	data_out_8,
	data_out_9,
	reset_n,
	clr_break_line,
	d_write,
	mem_used_1,
	Equal4,
	wait_latency_counter_1,
	wait_latency_counter_0,
	M_alu_result_3,
	M_alu_result_2,
	readdata_0,
	readdata_8,
	readdata_5,
	readdata_4,
	readdata_6,
	readdata_7,
	readdata_9,
	readdata_3,
	readdata_2,
	readdata_1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	[31:0] writedata;
output 	data_out_0;
output 	data_out_1;
output 	data_out_2;
output 	data_out_3;
output 	data_out_4;
output 	data_out_5;
output 	data_out_6;
output 	data_out_7;
output 	data_out_8;
output 	data_out_9;
input 	reset_n;
input 	clr_break_line;
input 	d_write;
input 	mem_used_1;
input 	Equal4;
input 	wait_latency_counter_1;
input 	wait_latency_counter_0;
input 	M_alu_result_3;
input 	M_alu_result_2;
output 	readdata_0;
output 	readdata_8;
output 	readdata_5;
output 	readdata_4;
output 	readdata_6;
output 	readdata_7;
output 	readdata_9;
output 	readdata_3;
output 	readdata_2;
output 	readdata_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \always0~0_combout ;
wire \always0~1_combout ;


dffeas \data_out[0] (
	.clk(clk),
	.d(writedata[0]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(data_out_0),
	.prn(vcc));
defparam \data_out[0] .is_wysiwyg = "true";
defparam \data_out[0] .power_up = "low";

dffeas \data_out[1] (
	.clk(clk),
	.d(writedata[1]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(data_out_1),
	.prn(vcc));
defparam \data_out[1] .is_wysiwyg = "true";
defparam \data_out[1] .power_up = "low";

dffeas \data_out[2] (
	.clk(clk),
	.d(writedata[2]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(data_out_2),
	.prn(vcc));
defparam \data_out[2] .is_wysiwyg = "true";
defparam \data_out[2] .power_up = "low";

dffeas \data_out[3] (
	.clk(clk),
	.d(writedata[3]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(data_out_3),
	.prn(vcc));
defparam \data_out[3] .is_wysiwyg = "true";
defparam \data_out[3] .power_up = "low";

dffeas \data_out[4] (
	.clk(clk),
	.d(writedata[4]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(data_out_4),
	.prn(vcc));
defparam \data_out[4] .is_wysiwyg = "true";
defparam \data_out[4] .power_up = "low";

dffeas \data_out[5] (
	.clk(clk),
	.d(writedata[5]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(data_out_5),
	.prn(vcc));
defparam \data_out[5] .is_wysiwyg = "true";
defparam \data_out[5] .power_up = "low";

dffeas \data_out[6] (
	.clk(clk),
	.d(writedata[6]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(data_out_6),
	.prn(vcc));
defparam \data_out[6] .is_wysiwyg = "true";
defparam \data_out[6] .power_up = "low";

dffeas \data_out[7] (
	.clk(clk),
	.d(writedata[7]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(data_out_7),
	.prn(vcc));
defparam \data_out[7] .is_wysiwyg = "true";
defparam \data_out[7] .power_up = "low";

dffeas \data_out[8] (
	.clk(clk),
	.d(writedata[8]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(data_out_8),
	.prn(vcc));
defparam \data_out[8] .is_wysiwyg = "true";
defparam \data_out[8] .power_up = "low";

dffeas \data_out[9] (
	.clk(clk),
	.d(writedata[9]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(data_out_9),
	.prn(vcc));
defparam \data_out[9] .is_wysiwyg = "true";
defparam \data_out[9] .power_up = "low";

cyclonev_lcell_comb \readdata[0] (
	.dataa(!data_out_0),
	.datab(!M_alu_result_3),
	.datac(!M_alu_result_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(readdata_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata[0] .extended_lut = "off";
defparam \readdata[0] .lut_mask = 64'hFDFDFDFDFDFDFDFD;
defparam \readdata[0] .shared_arith = "off";

cyclonev_lcell_comb \readdata[8] (
	.dataa(!data_out_8),
	.datab(!M_alu_result_3),
	.datac(!M_alu_result_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(readdata_8),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata[8] .extended_lut = "off";
defparam \readdata[8] .lut_mask = 64'hFDFDFDFDFDFDFDFD;
defparam \readdata[8] .shared_arith = "off";

cyclonev_lcell_comb \readdata[5] (
	.dataa(!data_out_5),
	.datab(!M_alu_result_3),
	.datac(!M_alu_result_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(readdata_5),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata[5] .extended_lut = "off";
defparam \readdata[5] .lut_mask = 64'hFDFDFDFDFDFDFDFD;
defparam \readdata[5] .shared_arith = "off";

cyclonev_lcell_comb \readdata[4] (
	.dataa(!data_out_4),
	.datab(!M_alu_result_3),
	.datac(!M_alu_result_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(readdata_4),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata[4] .extended_lut = "off";
defparam \readdata[4] .lut_mask = 64'hFDFDFDFDFDFDFDFD;
defparam \readdata[4] .shared_arith = "off";

cyclonev_lcell_comb \readdata[6] (
	.dataa(!data_out_6),
	.datab(!M_alu_result_3),
	.datac(!M_alu_result_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(readdata_6),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata[6] .extended_lut = "off";
defparam \readdata[6] .lut_mask = 64'hFDFDFDFDFDFDFDFD;
defparam \readdata[6] .shared_arith = "off";

cyclonev_lcell_comb \readdata[7] (
	.dataa(!data_out_7),
	.datab(!M_alu_result_3),
	.datac(!M_alu_result_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(readdata_7),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata[7] .extended_lut = "off";
defparam \readdata[7] .lut_mask = 64'hFDFDFDFDFDFDFDFD;
defparam \readdata[7] .shared_arith = "off";

cyclonev_lcell_comb \readdata[9] (
	.dataa(!data_out_9),
	.datab(!M_alu_result_3),
	.datac(!M_alu_result_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(readdata_9),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata[9] .extended_lut = "off";
defparam \readdata[9] .lut_mask = 64'hFDFDFDFDFDFDFDFD;
defparam \readdata[9] .shared_arith = "off";

cyclonev_lcell_comb \readdata[3] (
	.dataa(!data_out_3),
	.datab(!M_alu_result_3),
	.datac(!M_alu_result_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(readdata_3),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata[3] .extended_lut = "off";
defparam \readdata[3] .lut_mask = 64'hFDFDFDFDFDFDFDFD;
defparam \readdata[3] .shared_arith = "off";

cyclonev_lcell_comb \readdata[2] (
	.dataa(!data_out_2),
	.datab(!M_alu_result_3),
	.datac(!M_alu_result_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(readdata_2),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata[2] .extended_lut = "off";
defparam \readdata[2] .lut_mask = 64'hFDFDFDFDFDFDFDFD;
defparam \readdata[2] .shared_arith = "off";

cyclonev_lcell_comb \readdata[1] (
	.dataa(!data_out_1),
	.datab(!M_alu_result_3),
	.datac(!M_alu_result_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(readdata_1),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata[1] .extended_lut = "off";
defparam \readdata[1] .lut_mask = 64'hFDFDFDFDFDFDFDFD;
defparam \readdata[1] .shared_arith = "off";

cyclonev_lcell_comb \always0~0 (
	.dataa(!wait_latency_counter_1),
	.datab(!wait_latency_counter_0),
	.datac(!M_alu_result_3),
	.datad(!M_alu_result_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always0~0 .extended_lut = "off";
defparam \always0~0 .lut_mask = 64'hFFFEFFFEFFFEFFFE;
defparam \always0~0 .shared_arith = "off";

cyclonev_lcell_comb \always0~1 (
	.dataa(!clr_break_line),
	.datab(!d_write),
	.datac(!mem_used_1),
	.datad(!Equal4),
	.datae(!\always0~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always0~1 .extended_lut = "off";
defparam \always0~1 .lut_mask = 64'hF7FFFFFFF7FFFFFF;
defparam \always0~1 .shared_arith = "off";

endmodule

module processor_processor_mm_interconnect_0 (
	M_st_data_8,
	M_st_data_9,
	q_a_0,
	q_a_16,
	q_a_8,
	q_a_24,
	q_a_5,
	q_a_21,
	q_a_13,
	q_a_29,
	q_a_4,
	q_a_20,
	q_a_12,
	q_a_28,
	q_a_6,
	q_a_22,
	q_a_14,
	q_a_30,
	q_a_7,
	q_a_23,
	q_a_15,
	q_a_31,
	q_a_11,
	q_a_27,
	q_a_10,
	q_a_26,
	q_a_25,
	q_a_9,
	q_a_3,
	q_a_19,
	q_a_2,
	q_a_18,
	q_a_1,
	q_a_17,
	readdata_0,
	q_b_0,
	Add1,
	readdata_16,
	M_st_data_16,
	readdata_8,
	readdata_24,
	readdata_5,
	q_b_5,
	readdata_21,
	M_st_data_21,
	Add11,
	readdata_13,
	M_st_data_13,
	readdata_29,
	readdata_4,
	q_b_4,
	readdata_20,
	M_st_data_20,
	Add12,
	readdata_12,
	M_st_data_12,
	readdata_28,
	readdata_6,
	q_b_6,
	readdata_22,
	M_st_data_22,
	Add13,
	readdata_14,
	M_st_data_14,
	readdata_30,
	readdata_7,
	q_b_7,
	readdata_23,
	M_st_data_23,
	readdata_15,
	M_st_data_15,
	readdata_31,
	readdata_11,
	M_st_data_11,
	readdata_27,
	readdata_10,
	M_st_data_10,
	readdata_26,
	readdata_25,
	readdata_9,
	q_b_3,
	readdata_3,
	readdata_19,
	M_st_data_19,
	Add14,
	q_b_2,
	readdata_2,
	Add15,
	readdata_18,
	M_st_data_18,
	q_b_1,
	readdata_1,
	readdata_17,
	M_st_data_17,
	Add16,
	M_st_data_0,
	r_sync_rst,
	clr_break_line,
	d_write,
	mem_used_1,
	M_alu_result_5,
	M_alu_result_4,
	M_alu_result_6,
	M_alu_result_16,
	M_alu_result_15,
	M_alu_result_14,
	M_alu_result_13,
	Equal1,
	M_alu_result_12,
	M_alu_result_11,
	M_alu_result_10,
	M_alu_result_9,
	M_alu_result_8,
	M_alu_result_7,
	Equal2,
	Equal4,
	wait_latency_counter_1,
	wait_latency_counter_0,
	M_alu_result_3,
	M_alu_result_2,
	M_st_data_1,
	M_st_data_2,
	M_st_data_3,
	M_st_data_4,
	M_st_data_5,
	M_st_data_6,
	M_st_data_7,
	d_read,
	WideOr1,
	read_accepted,
	mem_used_11,
	wait_latency_counter_11,
	wait_latency_counter_01,
	av_waitrequest,
	Equal6,
	saved_grant_0,
	waitrequest,
	mem_used_12,
	saved_grant_01,
	mem_used_13,
	read_accepted1,
	hbreak_enabled,
	uav_read,
	src2_valid,
	saved_grant_1,
	i_read,
	has_pending_responses,
	ic_fill_tag_5,
	ic_fill_tag_4,
	ic_fill_tag_3,
	ic_fill_tag_2,
	ic_fill_tag_1,
	ic_fill_tag_0,
	Equal11,
	src0_valid,
	rf_source_valid,
	src3_valid,
	saved_grant_11,
	last_dest_id_1,
	src1_valid,
	read_latency_shift_reg,
	period_l_wr_strobe,
	src_data_0,
	src_payload,
	src_data_8,
	src_payload1,
	WideOr0,
	nonposted_cmd_accepted,
	ic_fill_line_5,
	src_data_46,
	src_data_5,
	src_payload2,
	src_payload3,
	src_payload4,
	src_data_4,
	src_payload5,
	src_payload6,
	src_payload7,
	src_data_6,
	src_payload8,
	src_payload9,
	src_payload10,
	src_data_7,
	src_payload11,
	src_payload12,
	src_payload13,
	ien_AE,
	av_readdata_9,
	ien_AF,
	av_readdata_8,
	src_payload14,
	src_payload15,
	src_payload16,
	src_payload17,
	src_payload18,
	src_data_9,
	src_data_3,
	src_payload19,
	src_data_2,
	src_payload20,
	src_data_1,
	src_payload21,
	b_full,
	ic_fill_line_0,
	ic_fill_line_1,
	ic_fill_line_2,
	ic_fill_line_3,
	ic_fill_line_4,
	src_payload22,
	ic_fill_ap_offset_0,
	src_data_38,
	ic_fill_ap_offset_1,
	src_data_39,
	ic_fill_ap_offset_2,
	src_data_40,
	src_data_41,
	src_data_42,
	src_data_43,
	src_data_44,
	src_data_45,
	src_data_461,
	src_data_47,
	src_data_48,
	src_data_49,
	src_data_50,
	M_mem_byte_en_0,
	src_data_32,
	readdata_01,
	readdata_02,
	read_0,
	readdata_03,
	counter_reg_bit_0,
	src_payload23,
	M_mem_byte_en_2,
	src_data_34,
	src_payload24,
	M_mem_byte_en_1,
	src_data_33,
	readdata_81,
	readdata_82,
	readdata_83,
	M_st_data_24,
	src_payload25,
	M_mem_byte_en_3,
	src_data_35,
	src_payload26,
	src_data_381,
	src_data_411,
	src_data_401,
	src_data_391,
	src_data_451,
	src_data_441,
	src_data_431,
	src_data_421,
	src_payload27,
	src_payload28,
	readdata_51,
	readdata_52,
	readdata_53,
	src_payload29,
	counter_reg_bit_5,
	src_payload30,
	b_full1,
	readdata_131,
	M_st_data_29,
	src_payload31,
	src_payload32,
	readdata_41,
	readdata_42,
	readdata_43,
	src_payload33,
	counter_reg_bit_4,
	src_payload34,
	b_non_empty,
	readdata_121,
	M_st_data_28,
	src_payload35,
	src_payload36,
	readdata_61,
	readdata_62,
	readdata_63,
	src_payload37,
	src_payload38,
	woverflow,
	readdata_141,
	M_st_data_30,
	src_payload39,
	src_payload40,
	readdata_71,
	readdata_72,
	readdata_73,
	src_payload41,
	src_payload42,
	rvalid,
	readdata_151,
	M_st_data_31,
	src_payload43,
	src_payload44,
	readdata_111,
	M_st_data_27,
	src_payload45,
	src_payload46,
	ac,
	readdata_101,
	M_st_data_26,
	src_payload47,
	M_st_data_25,
	src_payload48,
	src_payload49,
	readdata_91,
	readdata_92,
	readdata_93,
	src_payload50,
	readdata_32,
	readdata_33,
	readdata_34,
	src_payload51,
	counter_reg_bit_3,
	src_payload52,
	readdata_210,
	readdata_211,
	readdata_212,
	counter_reg_bit_2,
	src_payload53,
	src_payload54,
	readdata_110,
	readdata_112,
	readdata_113,
	src_payload55,
	counter_reg_bit_1,
	src_payload56,
	src_data_321,
	WideOr11,
	src_data_24,
	src_data_01,
	src_data_11,
	src_data_21,
	src_data_31,
	src_data_410,
	src_data_51,
	src_data_22,
	src_data_23,
	src_data_25,
	src_data_26,
	src_data_14,
	src_data_12,
	src_data_111,
	src_data_16,
	src_data_15,
	src_data_13,
	src_data_211,
	src_data_29,
	src_data_27,
	src_data_28,
	src_data_30,
	src_data_311,
	src_data_10,
	src_data_61,
	src_data_81,
	src_payload57,
	src_data_71,
	src_data_20,
	src_data_19,
	src_data_18,
	src_data_17,
	src_data_91,
	src_payload58,
	src_payload59,
	src_data_341,
	src_payload60,
	src_data_331,
	src_payload61,
	src_data_351,
	src_payload62,
	src_payload63,
	src_payload64,
	src_payload65,
	src_payload66,
	src_payload67,
	src_payload68,
	src_payload69,
	src_payload70,
	src_payload71,
	src_payload72,
	src_payload73,
	src_payload74,
	src_payload75,
	src_payload76,
	src_payload77,
	src_payload78,
	src_payload79,
	src_payload80,
	src_payload81,
	src_payload82,
	src_payload83,
	src_payload84,
	src_payload85,
	src_payload86,
	GND_port,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	M_st_data_8;
input 	M_st_data_9;
input 	q_a_0;
input 	q_a_16;
input 	q_a_8;
input 	q_a_24;
input 	q_a_5;
input 	q_a_21;
input 	q_a_13;
input 	q_a_29;
input 	q_a_4;
input 	q_a_20;
input 	q_a_12;
input 	q_a_28;
input 	q_a_6;
input 	q_a_22;
input 	q_a_14;
input 	q_a_30;
input 	q_a_7;
input 	q_a_23;
input 	q_a_15;
input 	q_a_31;
input 	q_a_11;
input 	q_a_27;
input 	q_a_10;
input 	q_a_26;
input 	q_a_25;
input 	q_a_9;
input 	q_a_3;
input 	q_a_19;
input 	q_a_2;
input 	q_a_18;
input 	q_a_1;
input 	q_a_17;
input 	readdata_0;
input 	q_b_0;
input 	Add1;
input 	readdata_16;
input 	M_st_data_16;
input 	readdata_8;
input 	readdata_24;
input 	readdata_5;
input 	q_b_5;
input 	readdata_21;
input 	M_st_data_21;
input 	Add11;
input 	readdata_13;
input 	M_st_data_13;
input 	readdata_29;
input 	readdata_4;
input 	q_b_4;
input 	readdata_20;
input 	M_st_data_20;
input 	Add12;
input 	readdata_12;
input 	M_st_data_12;
input 	readdata_28;
input 	readdata_6;
input 	q_b_6;
input 	readdata_22;
input 	M_st_data_22;
input 	Add13;
input 	readdata_14;
input 	M_st_data_14;
input 	readdata_30;
input 	readdata_7;
input 	q_b_7;
input 	readdata_23;
input 	M_st_data_23;
input 	readdata_15;
input 	M_st_data_15;
input 	readdata_31;
input 	readdata_11;
input 	M_st_data_11;
input 	readdata_27;
input 	readdata_10;
input 	M_st_data_10;
input 	readdata_26;
input 	readdata_25;
input 	readdata_9;
input 	q_b_3;
input 	readdata_3;
input 	readdata_19;
input 	M_st_data_19;
input 	Add14;
input 	q_b_2;
input 	readdata_2;
input 	Add15;
input 	readdata_18;
input 	M_st_data_18;
input 	q_b_1;
input 	readdata_1;
input 	readdata_17;
input 	M_st_data_17;
input 	Add16;
input 	M_st_data_0;
input 	r_sync_rst;
input 	clr_break_line;
input 	d_write;
output 	mem_used_1;
input 	M_alu_result_5;
input 	M_alu_result_4;
input 	M_alu_result_6;
input 	M_alu_result_16;
input 	M_alu_result_15;
input 	M_alu_result_14;
input 	M_alu_result_13;
output 	Equal1;
input 	M_alu_result_12;
input 	M_alu_result_11;
input 	M_alu_result_10;
input 	M_alu_result_9;
input 	M_alu_result_8;
input 	M_alu_result_7;
output 	Equal2;
output 	Equal4;
output 	wait_latency_counter_1;
output 	wait_latency_counter_0;
input 	M_alu_result_3;
input 	M_alu_result_2;
input 	M_st_data_1;
input 	M_st_data_2;
input 	M_st_data_3;
input 	M_st_data_4;
input 	M_st_data_5;
input 	M_st_data_6;
input 	M_st_data_7;
input 	d_read;
output 	WideOr1;
output 	read_accepted;
output 	mem_used_11;
output 	wait_latency_counter_11;
output 	wait_latency_counter_01;
input 	av_waitrequest;
output 	Equal6;
output 	saved_grant_0;
input 	waitrequest;
output 	mem_used_12;
output 	saved_grant_01;
output 	mem_used_13;
output 	read_accepted1;
input 	hbreak_enabled;
output 	uav_read;
output 	src2_valid;
output 	saved_grant_1;
input 	i_read;
output 	has_pending_responses;
input 	ic_fill_tag_5;
input 	ic_fill_tag_4;
input 	ic_fill_tag_3;
input 	ic_fill_tag_2;
input 	ic_fill_tag_1;
input 	ic_fill_tag_0;
output 	Equal11;
output 	src0_valid;
output 	rf_source_valid;
output 	src3_valid;
output 	saved_grant_11;
output 	last_dest_id_1;
output 	src1_valid;
output 	read_latency_shift_reg;
input 	period_l_wr_strobe;
output 	src_data_0;
output 	src_payload;
output 	src_data_8;
output 	src_payload1;
output 	WideOr0;
output 	nonposted_cmd_accepted;
input 	ic_fill_line_5;
output 	src_data_46;
output 	src_data_5;
output 	src_payload2;
output 	src_payload3;
output 	src_payload4;
output 	src_data_4;
output 	src_payload5;
output 	src_payload6;
output 	src_payload7;
output 	src_data_6;
output 	src_payload8;
output 	src_payload9;
output 	src_payload10;
output 	src_data_7;
output 	src_payload11;
output 	src_payload12;
output 	src_payload13;
input 	ien_AE;
input 	av_readdata_9;
input 	ien_AF;
input 	av_readdata_8;
output 	src_payload14;
output 	src_payload15;
output 	src_payload16;
output 	src_payload17;
output 	src_payload18;
output 	src_data_9;
output 	src_data_3;
output 	src_payload19;
output 	src_data_2;
output 	src_payload20;
output 	src_data_1;
output 	src_payload21;
input 	b_full;
input 	ic_fill_line_0;
input 	ic_fill_line_1;
input 	ic_fill_line_2;
input 	ic_fill_line_3;
input 	ic_fill_line_4;
output 	src_payload22;
input 	ic_fill_ap_offset_0;
output 	src_data_38;
input 	ic_fill_ap_offset_1;
output 	src_data_39;
input 	ic_fill_ap_offset_2;
output 	src_data_40;
output 	src_data_41;
output 	src_data_42;
output 	src_data_43;
output 	src_data_44;
output 	src_data_45;
output 	src_data_461;
output 	src_data_47;
output 	src_data_48;
output 	src_data_49;
output 	src_data_50;
input 	M_mem_byte_en_0;
output 	src_data_32;
input 	readdata_01;
input 	readdata_02;
input 	read_0;
input 	readdata_03;
input 	counter_reg_bit_0;
output 	src_payload23;
input 	M_mem_byte_en_2;
output 	src_data_34;
output 	src_payload24;
input 	M_mem_byte_en_1;
output 	src_data_33;
input 	readdata_81;
input 	readdata_82;
input 	readdata_83;
input 	M_st_data_24;
output 	src_payload25;
input 	M_mem_byte_en_3;
output 	src_data_35;
output 	src_payload26;
output 	src_data_381;
output 	src_data_411;
output 	src_data_401;
output 	src_data_391;
output 	src_data_451;
output 	src_data_441;
output 	src_data_431;
output 	src_data_421;
output 	src_payload27;
output 	src_payload28;
input 	readdata_51;
input 	readdata_52;
input 	readdata_53;
output 	src_payload29;
input 	counter_reg_bit_5;
output 	src_payload30;
input 	b_full1;
input 	readdata_131;
input 	M_st_data_29;
output 	src_payload31;
output 	src_payload32;
input 	readdata_41;
input 	readdata_42;
input 	readdata_43;
output 	src_payload33;
input 	counter_reg_bit_4;
output 	src_payload34;
input 	b_non_empty;
input 	readdata_121;
input 	M_st_data_28;
output 	src_payload35;
output 	src_payload36;
input 	readdata_61;
input 	readdata_62;
input 	readdata_63;
output 	src_payload37;
output 	src_payload38;
input 	woverflow;
input 	readdata_141;
input 	M_st_data_30;
output 	src_payload39;
output 	src_payload40;
input 	readdata_71;
input 	readdata_72;
input 	readdata_73;
output 	src_payload41;
output 	src_payload42;
input 	rvalid;
input 	readdata_151;
input 	M_st_data_31;
output 	src_payload43;
output 	src_payload44;
input 	readdata_111;
input 	M_st_data_27;
output 	src_payload45;
output 	src_payload46;
input 	ac;
input 	readdata_101;
input 	M_st_data_26;
output 	src_payload47;
input 	M_st_data_25;
output 	src_payload48;
output 	src_payload49;
input 	readdata_91;
input 	readdata_92;
input 	readdata_93;
output 	src_payload50;
input 	readdata_32;
input 	readdata_33;
input 	readdata_34;
output 	src_payload51;
input 	counter_reg_bit_3;
output 	src_payload52;
input 	readdata_210;
input 	readdata_211;
input 	readdata_212;
input 	counter_reg_bit_2;
output 	src_payload53;
output 	src_payload54;
input 	readdata_110;
input 	readdata_112;
input 	readdata_113;
output 	src_payload55;
input 	counter_reg_bit_1;
output 	src_payload56;
output 	src_data_321;
output 	WideOr11;
output 	src_data_24;
output 	src_data_01;
output 	src_data_11;
output 	src_data_21;
output 	src_data_31;
output 	src_data_410;
output 	src_data_51;
output 	src_data_22;
output 	src_data_23;
output 	src_data_25;
output 	src_data_26;
output 	src_data_14;
output 	src_data_12;
output 	src_data_111;
output 	src_data_16;
output 	src_data_15;
output 	src_data_13;
output 	src_data_211;
output 	src_data_29;
output 	src_data_27;
output 	src_data_28;
output 	src_data_30;
output 	src_data_311;
output 	src_data_10;
output 	src_data_61;
output 	src_data_81;
output 	src_payload57;
output 	src_data_71;
output 	src_data_20;
output 	src_data_19;
output 	src_data_18;
output 	src_data_17;
output 	src_data_91;
output 	src_payload58;
output 	src_payload59;
output 	src_data_341;
output 	src_payload60;
output 	src_data_331;
output 	src_payload61;
output 	src_data_351;
output 	src_payload62;
output 	src_payload63;
output 	src_payload64;
output 	src_payload65;
output 	src_payload66;
output 	src_payload67;
output 	src_payload68;
output 	src_payload69;
output 	src_payload70;
output 	src_payload71;
output 	src_payload72;
output 	src_payload73;
output 	src_payload74;
output 	src_payload75;
output 	src_payload76;
output 	src_payload77;
output 	src_payload78;
output 	src_payload79;
output 	src_payload80;
output 	src_payload81;
output 	src_payload82;
output 	src_payload83;
output 	src_payload84;
output 	src_payload85;
output 	src_payload86;
input 	GND_port;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[0]~q ;
wire \jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[16]~q ;
wire \jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[5]~q ;
wire \jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[21]~q ;
wire \jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[4]~q ;
wire \jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[20]~q ;
wire \jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[6]~q ;
wire \jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[22]~q ;
wire \jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[7]~q ;
wire \jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[3]~q ;
wire \jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[19]~q ;
wire \jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[2]~q ;
wire \jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[18]~q ;
wire \jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[1]~q ;
wire \jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[17]~q ;
wire \switches_pio_s1_translator|read_latency_shift_reg[0]~q ;
wire \cpu_jtag_debug_module_translator|read_latency_shift_reg[0]~q ;
wire \cpu_jtag_debug_module_agent_rsp_fifo|mem[0][74]~q ;
wire \cpu_jtag_debug_module_agent_rsp_fifo|mem[0][56]~q ;
wire \rsp_demux_002|src0_valid~0_combout ;
wire \onchip_mem_s1_translator|read_latency_shift_reg[0]~q ;
wire \onchip_mem_s1_agent_rsp_fifo|mem[0][74]~q ;
wire \onchip_mem_s1_agent_rsp_fifo|mem[0][56]~q ;
wire \rsp_demux_003|src0_valid~0_combout ;
wire \jtag_uart_avalon_jtag_slave_translator|read_latency_shift_reg[0]~q ;
wire \sysid_control_slave_translator|read_latency_shift_reg[0]~q ;
wire \sys_clk_timer_s1_translator|read_latency_shift_reg[0]~q ;
wire \led_pio_s1_translator|read_latency_shift_reg[0]~q ;
wire \sysid_control_slave_agent_rsp_fifo|mem_used[1]~q ;
wire \router|always1~0_combout ;
wire \router|always1~1_combout ;
wire \cmd_demux|sink_ready~0_combout ;
wire \sysid_control_slave_translator|wait_latency_counter[1]~q ;
wire \sysid_control_slave_translator|wait_latency_counter[0]~q ;
wire \cmd_demux|sink_ready~1_combout ;
wire \switches_pio_s1_agent_rsp_fifo|mem_used[1]~q ;
wire \router|always1~2_combout ;
wire \cmd_demux|sink_ready~2_combout ;
wire \switches_pio_s1_translator|wait_latency_counter[1]~q ;
wire \switches_pio_s1_translator|wait_latency_counter[0]~q ;
wire \cmd_demux|sink_ready~3_combout ;
wire \router|Equal2~1_combout ;
wire \jtag_uart_avalon_jtag_slave_agent_rsp_fifo|mem_used[1]~q ;
wire \cmd_demux|sink_ready~4_combout ;
wire \cpu_jtag_debug_module_agent_rsp_fifo|write~0_combout ;
wire \onchip_mem_s1_translator|read_latency_shift_reg~0_combout ;
wire \router|Equal1~1_combout ;
wire \cmd_demux|WideOr0~0_combout ;
wire \cmd_demux|src2_valid~0_combout ;
wire \led_pio_s1_translator|av_waitrequest_generated~0_combout ;
wire \led_pio_s1_agent_rsp_fifo|mem_used[1]~0_combout ;
wire \cmd_demux|src2_valid~1_combout ;
wire \cpu_instruction_master_limiter|last_channel[0]~q ;
wire \onchip_mem_s1_agent|rf_source_valid~0_combout ;
wire \onchip_mem_s1_translator|read_latency_shift_reg~1_combout ;
wire \router|Equal6~1_combout ;
wire \sys_clk_timer_s1_agent_rsp_fifo|mem_used[1]~0_combout ;
wire \sys_clk_timer_s1_translator|read_latency_shift_reg~0_combout ;
wire \cmd_demux|sink_ready~5_combout ;
wire \cmd_demux|sink_ready~6_combout ;
wire \cmd_demux|sink_ready~7_combout ;
wire \cmd_demux|sink_ready~8_combout ;
wire \switches_pio_s1_translator|av_readdata_pre[0]~q ;
wire \cpu_jtag_debug_module_translator|av_readdata_pre[0]~q ;
wire \led_pio_s1_translator|av_readdata_pre[0]~q ;
wire \sysid_control_slave_translator|av_readdata_pre[30]~q ;
wire \sys_clk_timer_s1_translator|av_readdata_pre[0]~q ;
wire \cpu_jtag_debug_module_translator|av_readdata_pre[16]~q ;
wire \led_pio_s1_translator|av_readdata_pre[8]~q ;
wire \jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[8]~q ;
wire \sys_clk_timer_s1_translator|av_readdata_pre[8]~q ;
wire \cpu_jtag_debug_module_translator|av_readdata_pre[8]~q ;
wire \switches_pio_s1_translator|av_readdata_pre[8]~q ;
wire \cpu_jtag_debug_module_translator|av_readdata_pre[24]~q ;
wire \rsp_demux_002|src1_valid~0_combout ;
wire \rsp_demux_003|src1_valid~0_combout ;
wire \cpu_jtag_debug_module_agent_rsp_fifo|mem[0][61]~q ;
wire \onchip_mem_s1_agent_rsp_fifo|mem[0][61]~q ;
wire \switches_pio_s1_translator|av_readdata_pre[5]~q ;
wire \cpu_jtag_debug_module_translator|av_readdata_pre[5]~q ;
wire \led_pio_s1_translator|av_readdata_pre[5]~q ;
wire \sys_clk_timer_s1_translator|av_readdata_pre[5]~q ;
wire \cpu_jtag_debug_module_translator|av_readdata_pre[21]~q ;
wire \cpu_jtag_debug_module_translator|av_readdata_pre[13]~q ;
wire \jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[13]~q ;
wire \sys_clk_timer_s1_translator|av_readdata_pre[13]~q ;
wire \cpu_jtag_debug_module_translator|av_readdata_pre[29]~q ;
wire \switches_pio_s1_translator|av_readdata_pre[4]~q ;
wire \cpu_jtag_debug_module_translator|av_readdata_pre[4]~q ;
wire \led_pio_s1_translator|av_readdata_pre[4]~q ;
wire \sys_clk_timer_s1_translator|av_readdata_pre[4]~q ;
wire \cpu_jtag_debug_module_translator|av_readdata_pre[20]~q ;
wire \cpu_jtag_debug_module_translator|av_readdata_pre[12]~q ;
wire \jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[12]~q ;
wire \sys_clk_timer_s1_translator|av_readdata_pre[12]~q ;
wire \cpu_jtag_debug_module_translator|av_readdata_pre[28]~q ;
wire \switches_pio_s1_translator|av_readdata_pre[6]~q ;
wire \cpu_jtag_debug_module_translator|av_readdata_pre[6]~q ;
wire \led_pio_s1_translator|av_readdata_pre[6]~q ;
wire \sys_clk_timer_s1_translator|av_readdata_pre[6]~q ;
wire \cpu_jtag_debug_module_translator|av_readdata_pre[22]~q ;
wire \cpu_jtag_debug_module_translator|av_readdata_pre[14]~q ;
wire \jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[14]~q ;
wire \sys_clk_timer_s1_translator|av_readdata_pre[14]~q ;
wire \cpu_jtag_debug_module_translator|av_readdata_pre[30]~q ;
wire \switches_pio_s1_translator|av_readdata_pre[7]~q ;
wire \cpu_jtag_debug_module_translator|av_readdata_pre[7]~q ;
wire \led_pio_s1_translator|av_readdata_pre[7]~q ;
wire \sys_clk_timer_s1_translator|av_readdata_pre[7]~q ;
wire \cpu_jtag_debug_module_translator|av_readdata_pre[23]~q ;
wire \cpu_jtag_debug_module_translator|av_readdata_pre[15]~q ;
wire \jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[15]~q ;
wire \sys_clk_timer_s1_translator|av_readdata_pre[15]~q ;
wire \cpu_jtag_debug_module_translator|av_readdata_pre[31]~q ;
wire \cpu_jtag_debug_module_translator|av_readdata_pre[11]~q ;
wire \sys_clk_timer_s1_translator|av_readdata_pre[11]~q ;
wire \cpu_jtag_debug_module_translator|av_readdata_pre[27]~q ;
wire \cpu_jtag_debug_module_translator|av_readdata_pre[10]~q ;
wire \jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[10]~q ;
wire \sys_clk_timer_s1_translator|av_readdata_pre[10]~q ;
wire \cpu_jtag_debug_module_translator|av_readdata_pre[26]~q ;
wire \cpu_jtag_debug_module_translator|av_readdata_pre[25]~q ;
wire \led_pio_s1_translator|av_readdata_pre[9]~q ;
wire \jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[9]~q ;
wire \sys_clk_timer_s1_translator|av_readdata_pre[9]~q ;
wire \cpu_jtag_debug_module_translator|av_readdata_pre[9]~q ;
wire \switches_pio_s1_translator|av_readdata_pre[9]~q ;
wire \led_pio_s1_translator|av_readdata_pre[3]~q ;
wire \sys_clk_timer_s1_translator|av_readdata_pre[3]~q ;
wire \cpu_jtag_debug_module_translator|av_readdata_pre[3]~q ;
wire \switches_pio_s1_translator|av_readdata_pre[3]~q ;
wire \cpu_jtag_debug_module_translator|av_readdata_pre[19]~q ;
wire \led_pio_s1_translator|av_readdata_pre[2]~q ;
wire \sys_clk_timer_s1_translator|av_readdata_pre[2]~q ;
wire \cpu_jtag_debug_module_translator|av_readdata_pre[2]~q ;
wire \switches_pio_s1_translator|av_readdata_pre[2]~q ;
wire \cpu_jtag_debug_module_translator|av_readdata_pre[18]~q ;
wire \led_pio_s1_translator|av_readdata_pre[1]~q ;
wire \sys_clk_timer_s1_translator|av_readdata_pre[1]~q ;
wire \cpu_jtag_debug_module_translator|av_readdata_pre[1]~q ;
wire \switches_pio_s1_translator|av_readdata_pre[1]~q ;
wire \cpu_jtag_debug_module_translator|av_readdata_pre[17]~q ;


processor_altera_merlin_slave_agent_3 onchip_mem_s1_agent(
	.saved_grant_0(saved_grant_01),
	.uav_read(uav_read),
	.i_read(i_read),
	.src3_valid(src3_valid),
	.saved_grant_1(saved_grant_11),
	.src1_valid(src1_valid),
	.rf_source_valid(\onchip_mem_s1_agent|rf_source_valid~0_combout ));

processor_altera_avalon_sc_fifo cpu_jtag_debug_module_agent_rsp_fifo(
	.reset(r_sync_rst),
	.read_latency_shift_reg_0(\cpu_jtag_debug_module_translator|read_latency_shift_reg[0]~q ),
	.mem_74_0(\cpu_jtag_debug_module_agent_rsp_fifo|mem[0][74]~q ),
	.mem_56_0(\cpu_jtag_debug_module_agent_rsp_fifo|mem[0][56]~q ),
	.saved_grant_0(saved_grant_0),
	.waitrequest(waitrequest),
	.mem_used_1(mem_used_12),
	.write(\cpu_jtag_debug_module_agent_rsp_fifo|write~0_combout ),
	.uav_read(uav_read),
	.saved_grant_1(saved_grant_1),
	.i_read(i_read),
	.rf_source_valid(rf_source_valid),
	.mem_61_0(\cpu_jtag_debug_module_agent_rsp_fifo|mem[0][61]~q ),
	.clk(clk_clk));

processor_altera_merlin_slave_agent cpu_jtag_debug_module_agent(
	.saved_grant_0(saved_grant_0),
	.uav_read(uav_read),
	.src2_valid(src2_valid),
	.saved_grant_1(saved_grant_1),
	.i_read(i_read),
	.src0_valid(src0_valid),
	.rf_source_valid(rf_source_valid));

processor_altera_avalon_sc_fifo_6 sysid_control_slave_agent_rsp_fifo(
	.reset(r_sync_rst),
	.read_latency_shift_reg_0(\sysid_control_slave_translator|read_latency_shift_reg[0]~q ),
	.mem_used_1(\sysid_control_slave_agent_rsp_fifo|mem_used[1]~q ),
	.sink_ready(\cmd_demux|sink_ready~1_combout ),
	.sink_ready1(\cmd_demux|sink_ready~5_combout ),
	.sink_ready2(\cmd_demux|sink_ready~6_combout ),
	.clk(clk_clk));

processor_altera_avalon_sc_fifo_1 jtag_uart_avalon_jtag_slave_agent_rsp_fifo(
	.reset(r_sync_rst),
	.clr_break_line(clr_break_line),
	.read_latency_shift_reg_0(\jtag_uart_avalon_jtag_slave_translator|read_latency_shift_reg[0]~q ),
	.mem_used_1(\jtag_uart_avalon_jtag_slave_agent_rsp_fifo|mem_used[1]~q ),
	.av_waitrequest(av_waitrequest),
	.uav_read(uav_read),
	.Equal6(\router|Equal6~1_combout ),
	.clk(clk_clk));

processor_altera_merlin_slave_translator_4 switches_pio_s1_translator(
	.reset(r_sync_rst),
	.d_write(d_write),
	.read_latency_shift_reg_0(\switches_pio_s1_translator|read_latency_shift_reg[0]~q ),
	.sink_ready(\cmd_demux|sink_ready~2_combout ),
	.wait_latency_counter_1(\switches_pio_s1_translator|wait_latency_counter[1]~q ),
	.wait_latency_counter_0(\switches_pio_s1_translator|wait_latency_counter[0]~q ),
	.sink_ready1(\cmd_demux|sink_ready~3_combout ),
	.uav_read(uav_read),
	.av_readdata_pre_0(\switches_pio_s1_translator|av_readdata_pre[0]~q ),
	.av_readdata_pre_8(\switches_pio_s1_translator|av_readdata_pre[8]~q ),
	.av_readdata_pre_5(\switches_pio_s1_translator|av_readdata_pre[5]~q ),
	.av_readdata_pre_4(\switches_pio_s1_translator|av_readdata_pre[4]~q ),
	.av_readdata_pre_6(\switches_pio_s1_translator|av_readdata_pre[6]~q ),
	.av_readdata_pre_7(\switches_pio_s1_translator|av_readdata_pre[7]~q ),
	.av_readdata_pre_9(\switches_pio_s1_translator|av_readdata_pre[9]~q ),
	.av_readdata_pre_3(\switches_pio_s1_translator|av_readdata_pre[3]~q ),
	.av_readdata_pre_2(\switches_pio_s1_translator|av_readdata_pre[2]~q ),
	.av_readdata_pre_1(\switches_pio_s1_translator|av_readdata_pre[1]~q ),
	.av_readdata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,readdata_93,readdata_83,readdata_71,readdata_61,readdata_51,readdata_41,readdata_34,readdata_212,readdata_113,readdata_01}),
	.clk(clk_clk));

processor_altera_merlin_slave_translator_2 led_pio_s1_translator(
	.reset(r_sync_rst),
	.clr_break_line(clr_break_line),
	.d_write(d_write),
	.mem_used_1(mem_used_1),
	.Equal4(Equal4),
	.wait_latency_counter_1(wait_latency_counter_1),
	.wait_latency_counter_0(wait_latency_counter_0),
	.read_latency_shift_reg_0(\led_pio_s1_translator|read_latency_shift_reg[0]~q ),
	.av_waitrequest_generated(\led_pio_s1_translator|av_waitrequest_generated~0_combout ),
	.mem_used_11(\led_pio_s1_agent_rsp_fifo|mem_used[1]~0_combout ),
	.src2_valid(\cmd_demux|src2_valid~1_combout ),
	.av_readdata_pre_0(\led_pio_s1_translator|av_readdata_pre[0]~q ),
	.av_readdata_pre_8(\led_pio_s1_translator|av_readdata_pre[8]~q ),
	.av_readdata_pre_5(\led_pio_s1_translator|av_readdata_pre[5]~q ),
	.av_readdata_pre_4(\led_pio_s1_translator|av_readdata_pre[4]~q ),
	.av_readdata_pre_6(\led_pio_s1_translator|av_readdata_pre[6]~q ),
	.av_readdata_pre_7(\led_pio_s1_translator|av_readdata_pre[7]~q ),
	.av_readdata_pre_9(\led_pio_s1_translator|av_readdata_pre[9]~q ),
	.av_readdata_pre_3(\led_pio_s1_translator|av_readdata_pre[3]~q ),
	.av_readdata_pre_2(\led_pio_s1_translator|av_readdata_pre[2]~q ),
	.av_readdata_pre_1(\led_pio_s1_translator|av_readdata_pre[1]~q ),
	.av_readdata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,readdata_91,readdata_81,readdata_72,readdata_62,readdata_52,readdata_42,readdata_32,readdata_210,readdata_110,readdata_02}),
	.clk(clk_clk));

processor_altera_merlin_slave_translator_5 sys_clk_timer_s1_translator(
	.reset(r_sync_rst),
	.d_write(d_write),
	.read_latency_shift_reg_0(\sys_clk_timer_s1_translator|read_latency_shift_reg[0]~q ),
	.wait_latency_counter_1(wait_latency_counter_11),
	.wait_latency_counter_0(wait_latency_counter_01),
	.uav_read(uav_read),
	.period_l_wr_strobe(period_l_wr_strobe),
	.mem_used_1(\sys_clk_timer_s1_agent_rsp_fifo|mem_used[1]~0_combout ),
	.read_latency_shift_reg(\sys_clk_timer_s1_translator|read_latency_shift_reg~0_combout ),
	.av_readdata_pre_0(\sys_clk_timer_s1_translator|av_readdata_pre[0]~q ),
	.av_readdata_pre_8(\sys_clk_timer_s1_translator|av_readdata_pre[8]~q ),
	.av_readdata_pre_5(\sys_clk_timer_s1_translator|av_readdata_pre[5]~q ),
	.av_readdata_pre_13(\sys_clk_timer_s1_translator|av_readdata_pre[13]~q ),
	.av_readdata_pre_4(\sys_clk_timer_s1_translator|av_readdata_pre[4]~q ),
	.av_readdata_pre_12(\sys_clk_timer_s1_translator|av_readdata_pre[12]~q ),
	.av_readdata_pre_6(\sys_clk_timer_s1_translator|av_readdata_pre[6]~q ),
	.av_readdata_pre_14(\sys_clk_timer_s1_translator|av_readdata_pre[14]~q ),
	.av_readdata_pre_7(\sys_clk_timer_s1_translator|av_readdata_pre[7]~q ),
	.av_readdata_pre_15(\sys_clk_timer_s1_translator|av_readdata_pre[15]~q ),
	.av_readdata_pre_11(\sys_clk_timer_s1_translator|av_readdata_pre[11]~q ),
	.av_readdata_pre_10(\sys_clk_timer_s1_translator|av_readdata_pre[10]~q ),
	.av_readdata_pre_9(\sys_clk_timer_s1_translator|av_readdata_pre[9]~q ),
	.av_readdata_pre_3(\sys_clk_timer_s1_translator|av_readdata_pre[3]~q ),
	.av_readdata_pre_2(\sys_clk_timer_s1_translator|av_readdata_pre[2]~q ),
	.av_readdata_pre_1(\sys_clk_timer_s1_translator|av_readdata_pre[1]~q ),
	.av_readdata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,readdata_151,readdata_141,readdata_131,readdata_121,readdata_111,readdata_101,readdata_92,readdata_82,readdata_73,readdata_63,readdata_53,readdata_43,readdata_33,readdata_211,readdata_112,readdata_03}),
	.clk(clk_clk));

processor_altera_merlin_slave_translator_3 onchip_mem_s1_translator(
	.reset(r_sync_rst),
	.clr_break_line(clr_break_line),
	.read_latency_shift_reg_0(\onchip_mem_s1_translator|read_latency_shift_reg[0]~q ),
	.mem_used_1(mem_used_13),
	.read_latency_shift_reg(\onchip_mem_s1_translator|read_latency_shift_reg~0_combout ),
	.rf_source_valid(\onchip_mem_s1_agent|rf_source_valid~0_combout ),
	.read_latency_shift_reg1(\onchip_mem_s1_translator|read_latency_shift_reg~1_combout ),
	.clk(clk_clk));

processor_altera_merlin_slave_translator cpu_jtag_debug_module_translator(
	.av_readdata({readdata_31,readdata_30,readdata_29,readdata_28,readdata_27,readdata_26,readdata_25,readdata_24,readdata_23,readdata_22,readdata_21,readdata_20,readdata_19,readdata_18,readdata_17,readdata_16,readdata_15,readdata_14,readdata_13,readdata_12,readdata_11,readdata_10,readdata_9,
readdata_8,readdata_7,readdata_6,readdata_5,readdata_4,readdata_3,readdata_2,readdata_1,readdata_0}),
	.reset(r_sync_rst),
	.clr_break_line(clr_break_line),
	.read_latency_shift_reg_0(\cpu_jtag_debug_module_translator|read_latency_shift_reg[0]~q ),
	.write(\cpu_jtag_debug_module_agent_rsp_fifo|write~0_combout ),
	.rf_source_valid(rf_source_valid),
	.av_readdata_pre_0(\cpu_jtag_debug_module_translator|av_readdata_pre[0]~q ),
	.av_readdata_pre_16(\cpu_jtag_debug_module_translator|av_readdata_pre[16]~q ),
	.av_readdata_pre_8(\cpu_jtag_debug_module_translator|av_readdata_pre[8]~q ),
	.av_readdata_pre_24(\cpu_jtag_debug_module_translator|av_readdata_pre[24]~q ),
	.av_readdata_pre_5(\cpu_jtag_debug_module_translator|av_readdata_pre[5]~q ),
	.av_readdata_pre_21(\cpu_jtag_debug_module_translator|av_readdata_pre[21]~q ),
	.av_readdata_pre_13(\cpu_jtag_debug_module_translator|av_readdata_pre[13]~q ),
	.av_readdata_pre_29(\cpu_jtag_debug_module_translator|av_readdata_pre[29]~q ),
	.av_readdata_pre_4(\cpu_jtag_debug_module_translator|av_readdata_pre[4]~q ),
	.av_readdata_pre_20(\cpu_jtag_debug_module_translator|av_readdata_pre[20]~q ),
	.av_readdata_pre_12(\cpu_jtag_debug_module_translator|av_readdata_pre[12]~q ),
	.av_readdata_pre_28(\cpu_jtag_debug_module_translator|av_readdata_pre[28]~q ),
	.av_readdata_pre_6(\cpu_jtag_debug_module_translator|av_readdata_pre[6]~q ),
	.av_readdata_pre_22(\cpu_jtag_debug_module_translator|av_readdata_pre[22]~q ),
	.av_readdata_pre_14(\cpu_jtag_debug_module_translator|av_readdata_pre[14]~q ),
	.av_readdata_pre_30(\cpu_jtag_debug_module_translator|av_readdata_pre[30]~q ),
	.av_readdata_pre_7(\cpu_jtag_debug_module_translator|av_readdata_pre[7]~q ),
	.av_readdata_pre_23(\cpu_jtag_debug_module_translator|av_readdata_pre[23]~q ),
	.av_readdata_pre_15(\cpu_jtag_debug_module_translator|av_readdata_pre[15]~q ),
	.av_readdata_pre_31(\cpu_jtag_debug_module_translator|av_readdata_pre[31]~q ),
	.av_readdata_pre_11(\cpu_jtag_debug_module_translator|av_readdata_pre[11]~q ),
	.av_readdata_pre_27(\cpu_jtag_debug_module_translator|av_readdata_pre[27]~q ),
	.av_readdata_pre_10(\cpu_jtag_debug_module_translator|av_readdata_pre[10]~q ),
	.av_readdata_pre_26(\cpu_jtag_debug_module_translator|av_readdata_pre[26]~q ),
	.av_readdata_pre_25(\cpu_jtag_debug_module_translator|av_readdata_pre[25]~q ),
	.av_readdata_pre_9(\cpu_jtag_debug_module_translator|av_readdata_pre[9]~q ),
	.av_readdata_pre_3(\cpu_jtag_debug_module_translator|av_readdata_pre[3]~q ),
	.av_readdata_pre_19(\cpu_jtag_debug_module_translator|av_readdata_pre[19]~q ),
	.av_readdata_pre_2(\cpu_jtag_debug_module_translator|av_readdata_pre[2]~q ),
	.av_readdata_pre_18(\cpu_jtag_debug_module_translator|av_readdata_pre[18]~q ),
	.av_readdata_pre_1(\cpu_jtag_debug_module_translator|av_readdata_pre[1]~q ),
	.av_readdata_pre_17(\cpu_jtag_debug_module_translator|av_readdata_pre[17]~q ),
	.clk(clk_clk));

processor_altera_merlin_slave_translator_6 sysid_control_slave_translator(
	.reset(r_sync_rst),
	.d_write(d_write),
	.av_readdata({gnd,M_alu_result_2,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.read_latency_shift_reg_0(\sysid_control_slave_translator|read_latency_shift_reg[0]~q ),
	.sink_ready(\cmd_demux|sink_ready~0_combout ),
	.wait_latency_counter_1(\sysid_control_slave_translator|wait_latency_counter[1]~q ),
	.wait_latency_counter_0(\sysid_control_slave_translator|wait_latency_counter[0]~q ),
	.sink_ready1(\cmd_demux|sink_ready~1_combout ),
	.uav_read(uav_read),
	.av_readdata_pre_30(\sysid_control_slave_translator|av_readdata_pre[30]~q ),
	.clk(clk_clk));

processor_altera_merlin_slave_translator_1 jtag_uart_avalon_jtag_slave_translator(
	.av_readdata_pre_0(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[0]~q ),
	.av_readdata_pre_16(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[16]~q ),
	.av_readdata_pre_5(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[5]~q ),
	.av_readdata_pre_21(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[21]~q ),
	.av_readdata_pre_4(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[4]~q ),
	.av_readdata_pre_20(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[20]~q ),
	.av_readdata_pre_6(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[6]~q ),
	.av_readdata_pre_22(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[22]~q ),
	.av_readdata_pre_7(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[7]~q ),
	.av_readdata_pre_3(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[3]~q ),
	.av_readdata_pre_19(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[19]~q ),
	.av_readdata_pre_2(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[2]~q ),
	.av_readdata_pre_18(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[18]~q ),
	.av_readdata_pre_1(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[1]~q ),
	.av_readdata_pre_17(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[17]~q ),
	.q_b_0(q_b_0),
	.av_readdata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,Add13,Add11,Add12,Add14,Add15,Add16,Add1,rvalid,woverflow,gnd,b_non_empty,gnd,ac,av_readdata_9,av_readdata_8,GND_port,GND_port,GND_port,GND_port,GND_port,GND_port,ien_AE,ien_AF}),
	.q_b_5(q_b_5),
	.q_b_4(q_b_4),
	.q_b_6(q_b_6),
	.q_b_7(q_b_7),
	.q_b_3(q_b_3),
	.q_b_2(q_b_2),
	.q_b_1(q_b_1),
	.reset(r_sync_rst),
	.clr_break_line(clr_break_line),
	.read_latency_shift_reg_0(\jtag_uart_avalon_jtag_slave_translator|read_latency_shift_reg[0]~q ),
	.mem_used_1(\jtag_uart_avalon_jtag_slave_agent_rsp_fifo|mem_used[1]~q ),
	.av_waitrequest(av_waitrequest),
	.uav_read(uav_read),
	.Equal6(\router|Equal6~1_combout ),
	.read_latency_shift_reg(read_latency_shift_reg),
	.av_readdata_pre_8(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[8]~q ),
	.av_readdata_pre_13(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[13]~q ),
	.av_readdata_pre_12(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[12]~q ),
	.av_readdata_pre_14(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[14]~q ),
	.av_readdata_pre_15(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[15]~q ),
	.av_readdata_pre_10(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[10]~q ),
	.av_readdata_pre_9(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[9]~q ),
	.b_full(b_full),
	.read_0(read_0),
	.counter_reg_bit_0(counter_reg_bit_0),
	.counter_reg_bit_5(counter_reg_bit_5),
	.b_full1(b_full1),
	.counter_reg_bit_4(counter_reg_bit_4),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_1(counter_reg_bit_1),
	.clk(clk_clk));

processor_altera_merlin_master_translator cpu_data_master_translator(
	.reset(r_sync_rst),
	.clr_break_line(clr_break_line),
	.d_write(d_write),
	.mem_used_1(mem_used_1),
	.Equal4(Equal4),
	.wait_latency_counter_1(wait_latency_counter_1),
	.wait_latency_counter_0(wait_latency_counter_0),
	.d_read(d_read),
	.WideOr1(WideOr1),
	.read_accepted1(read_accepted),
	.sink_ready(\cmd_demux|sink_ready~1_combout ),
	.sink_ready1(\cmd_demux|sink_ready~3_combout ),
	.Equal2(\router|Equal2~1_combout ),
	.mem_used_11(mem_used_11),
	.wait_latency_counter_11(wait_latency_counter_11),
	.wait_latency_counter_01(wait_latency_counter_01),
	.sink_ready2(\cmd_demux|sink_ready~4_combout ),
	.WideOr0(\cmd_demux|WideOr0~0_combout ),
	.src2_valid(\cmd_demux|src2_valid~0_combout ),
	.read_accepted2(read_accepted1),
	.uav_read(uav_read),
	.clk(clk_clk));

processor_processor_mm_interconnect_0_rsp_mux_001 rsp_mux_001(
	.q_a_0(q_a_0),
	.q_a_16(q_a_16),
	.q_a_8(q_a_8),
	.q_a_24(q_a_24),
	.q_a_5(q_a_5),
	.q_a_21(q_a_21),
	.q_a_13(q_a_13),
	.q_a_29(q_a_29),
	.q_a_4(q_a_4),
	.q_a_20(q_a_20),
	.q_a_12(q_a_12),
	.q_a_28(q_a_28),
	.q_a_6(q_a_6),
	.q_a_22(q_a_22),
	.q_a_14(q_a_14),
	.q_a_30(q_a_30),
	.q_a_7(q_a_7),
	.q_a_23(q_a_23),
	.q_a_15(q_a_15),
	.q_a_31(q_a_31),
	.q_a_11(q_a_11),
	.q_a_27(q_a_27),
	.q_a_10(q_a_10),
	.q_a_26(q_a_26),
	.q_a_25(q_a_25),
	.q_a_9(q_a_9),
	.q_a_3(q_a_3),
	.q_a_19(q_a_19),
	.q_a_2(q_a_2),
	.q_a_18(q_a_18),
	.q_a_1(q_a_1),
	.q_a_17(q_a_17),
	.av_readdata_pre_0(\cpu_jtag_debug_module_translator|av_readdata_pre[0]~q ),
	.av_readdata_pre_16(\cpu_jtag_debug_module_translator|av_readdata_pre[16]~q ),
	.av_readdata_pre_8(\cpu_jtag_debug_module_translator|av_readdata_pre[8]~q ),
	.av_readdata_pre_24(\cpu_jtag_debug_module_translator|av_readdata_pre[24]~q ),
	.src1_valid(\rsp_demux_002|src1_valid~0_combout ),
	.src1_valid1(\rsp_demux_003|src1_valid~0_combout ),
	.av_readdata_pre_5(\cpu_jtag_debug_module_translator|av_readdata_pre[5]~q ),
	.av_readdata_pre_21(\cpu_jtag_debug_module_translator|av_readdata_pre[21]~q ),
	.av_readdata_pre_13(\cpu_jtag_debug_module_translator|av_readdata_pre[13]~q ),
	.av_readdata_pre_29(\cpu_jtag_debug_module_translator|av_readdata_pre[29]~q ),
	.av_readdata_pre_4(\cpu_jtag_debug_module_translator|av_readdata_pre[4]~q ),
	.av_readdata_pre_20(\cpu_jtag_debug_module_translator|av_readdata_pre[20]~q ),
	.av_readdata_pre_12(\cpu_jtag_debug_module_translator|av_readdata_pre[12]~q ),
	.av_readdata_pre_28(\cpu_jtag_debug_module_translator|av_readdata_pre[28]~q ),
	.av_readdata_pre_6(\cpu_jtag_debug_module_translator|av_readdata_pre[6]~q ),
	.av_readdata_pre_22(\cpu_jtag_debug_module_translator|av_readdata_pre[22]~q ),
	.av_readdata_pre_14(\cpu_jtag_debug_module_translator|av_readdata_pre[14]~q ),
	.av_readdata_pre_30(\cpu_jtag_debug_module_translator|av_readdata_pre[30]~q ),
	.av_readdata_pre_7(\cpu_jtag_debug_module_translator|av_readdata_pre[7]~q ),
	.av_readdata_pre_23(\cpu_jtag_debug_module_translator|av_readdata_pre[23]~q ),
	.av_readdata_pre_15(\cpu_jtag_debug_module_translator|av_readdata_pre[15]~q ),
	.av_readdata_pre_31(\cpu_jtag_debug_module_translator|av_readdata_pre[31]~q ),
	.av_readdata_pre_11(\cpu_jtag_debug_module_translator|av_readdata_pre[11]~q ),
	.av_readdata_pre_27(\cpu_jtag_debug_module_translator|av_readdata_pre[27]~q ),
	.av_readdata_pre_10(\cpu_jtag_debug_module_translator|av_readdata_pre[10]~q ),
	.av_readdata_pre_26(\cpu_jtag_debug_module_translator|av_readdata_pre[26]~q ),
	.av_readdata_pre_25(\cpu_jtag_debug_module_translator|av_readdata_pre[25]~q ),
	.av_readdata_pre_9(\cpu_jtag_debug_module_translator|av_readdata_pre[9]~q ),
	.av_readdata_pre_3(\cpu_jtag_debug_module_translator|av_readdata_pre[3]~q ),
	.av_readdata_pre_19(\cpu_jtag_debug_module_translator|av_readdata_pre[19]~q ),
	.av_readdata_pre_2(\cpu_jtag_debug_module_translator|av_readdata_pre[2]~q ),
	.av_readdata_pre_18(\cpu_jtag_debug_module_translator|av_readdata_pre[18]~q ),
	.av_readdata_pre_1(\cpu_jtag_debug_module_translator|av_readdata_pre[1]~q ),
	.av_readdata_pre_17(\cpu_jtag_debug_module_translator|av_readdata_pre[17]~q ),
	.WideOr11(WideOr11),
	.src_data_24(src_data_24),
	.src_data_0(src_data_01),
	.src_data_1(src_data_11),
	.src_data_2(src_data_21),
	.src_data_3(src_data_31),
	.src_data_4(src_data_410),
	.src_data_5(src_data_51),
	.src_data_22(src_data_22),
	.src_data_23(src_data_23),
	.src_data_25(src_data_25),
	.src_data_26(src_data_26),
	.src_data_14(src_data_14),
	.src_data_12(src_data_12),
	.src_data_11(src_data_111),
	.src_data_16(src_data_16),
	.src_data_15(src_data_15),
	.src_data_13(src_data_13),
	.src_data_21(src_data_211),
	.src_data_29(src_data_29),
	.src_data_27(src_data_27),
	.src_data_28(src_data_28),
	.src_data_30(src_data_30),
	.src_data_31(src_data_311),
	.src_data_10(src_data_10),
	.src_data_6(src_data_61),
	.src_data_8(src_data_81),
	.src_data_7(src_data_71),
	.src_data_20(src_data_20),
	.src_data_19(src_data_19),
	.src_data_18(src_data_18),
	.src_data_17(src_data_17),
	.src_data_9(src_data_91));

processor_processor_mm_interconnect_0_rsp_mux rsp_mux(
	.q_a_0(q_a_0),
	.av_readdata_pre_0(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[0]~q ),
	.av_readdata_pre_16(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[16]~q ),
	.q_a_16(q_a_16),
	.q_a_8(q_a_8),
	.q_a_24(q_a_24),
	.q_a_5(q_a_5),
	.av_readdata_pre_5(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[5]~q ),
	.q_a_21(q_a_21),
	.av_readdata_pre_21(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[21]~q ),
	.q_a_13(q_a_13),
	.q_a_29(q_a_29),
	.q_a_4(q_a_4),
	.av_readdata_pre_4(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[4]~q ),
	.q_a_20(q_a_20),
	.av_readdata_pre_20(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[20]~q ),
	.q_a_12(q_a_12),
	.q_a_28(q_a_28),
	.q_a_6(q_a_6),
	.av_readdata_pre_6(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[6]~q ),
	.q_a_22(q_a_22),
	.av_readdata_pre_22(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[22]~q ),
	.q_a_14(q_a_14),
	.q_a_30(q_a_30),
	.q_a_7(q_a_7),
	.av_readdata_pre_7(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[7]~q ),
	.q_a_23(q_a_23),
	.q_a_15(q_a_15),
	.q_a_31(q_a_31),
	.q_a_11(q_a_11),
	.q_a_27(q_a_27),
	.q_a_10(q_a_10),
	.q_a_26(q_a_26),
	.q_a_25(q_a_25),
	.q_a_9(q_a_9),
	.q_a_3(q_a_3),
	.av_readdata_pre_3(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[3]~q ),
	.q_a_19(q_a_19),
	.av_readdata_pre_19(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[19]~q ),
	.q_a_2(q_a_2),
	.av_readdata_pre_2(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[2]~q ),
	.av_readdata_pre_18(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[18]~q ),
	.q_a_18(q_a_18),
	.q_a_1(q_a_1),
	.av_readdata_pre_1(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[1]~q ),
	.q_a_17(q_a_17),
	.av_readdata_pre_17(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[17]~q ),
	.read_latency_shift_reg_0(\switches_pio_s1_translator|read_latency_shift_reg[0]~q ),
	.src0_valid(\rsp_demux_002|src0_valid~0_combout ),
	.src0_valid1(\rsp_demux_003|src0_valid~0_combout ),
	.read_latency_shift_reg_01(\jtag_uart_avalon_jtag_slave_translator|read_latency_shift_reg[0]~q ),
	.read_latency_shift_reg_02(\sysid_control_slave_translator|read_latency_shift_reg[0]~q ),
	.read_latency_shift_reg_03(\sys_clk_timer_s1_translator|read_latency_shift_reg[0]~q ),
	.read_latency_shift_reg_04(\led_pio_s1_translator|read_latency_shift_reg[0]~q ),
	.WideOr11(WideOr1),
	.av_readdata_pre_01(\switches_pio_s1_translator|av_readdata_pre[0]~q ),
	.av_readdata_pre_02(\cpu_jtag_debug_module_translator|av_readdata_pre[0]~q ),
	.av_readdata_pre_03(\led_pio_s1_translator|av_readdata_pre[0]~q ),
	.av_readdata_pre_30(\sysid_control_slave_translator|av_readdata_pre[30]~q ),
	.av_readdata_pre_04(\sys_clk_timer_s1_translator|av_readdata_pre[0]~q ),
	.src_data_0(src_data_0),
	.av_readdata_pre_161(\cpu_jtag_debug_module_translator|av_readdata_pre[16]~q ),
	.src_payload(src_payload),
	.av_readdata_pre_8(\led_pio_s1_translator|av_readdata_pre[8]~q ),
	.av_readdata_pre_81(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[8]~q ),
	.av_readdata_pre_82(\sys_clk_timer_s1_translator|av_readdata_pre[8]~q ),
	.av_readdata_pre_83(\cpu_jtag_debug_module_translator|av_readdata_pre[8]~q ),
	.av_readdata_pre_84(\switches_pio_s1_translator|av_readdata_pre[8]~q ),
	.src_data_8(src_data_8),
	.av_readdata_pre_24(\cpu_jtag_debug_module_translator|av_readdata_pre[24]~q ),
	.src_payload1(src_payload1),
	.av_readdata_pre_51(\switches_pio_s1_translator|av_readdata_pre[5]~q ),
	.av_readdata_pre_52(\cpu_jtag_debug_module_translator|av_readdata_pre[5]~q ),
	.av_readdata_pre_53(\led_pio_s1_translator|av_readdata_pre[5]~q ),
	.av_readdata_pre_54(\sys_clk_timer_s1_translator|av_readdata_pre[5]~q ),
	.src_data_5(src_data_5),
	.av_readdata_pre_211(\cpu_jtag_debug_module_translator|av_readdata_pre[21]~q ),
	.src_payload2(src_payload2),
	.av_readdata_pre_13(\cpu_jtag_debug_module_translator|av_readdata_pre[13]~q ),
	.av_readdata_pre_131(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[13]~q ),
	.av_readdata_pre_132(\sys_clk_timer_s1_translator|av_readdata_pre[13]~q ),
	.src_payload3(src_payload3),
	.av_readdata_pre_29(\cpu_jtag_debug_module_translator|av_readdata_pre[29]~q ),
	.src_payload4(src_payload4),
	.av_readdata_pre_41(\switches_pio_s1_translator|av_readdata_pre[4]~q ),
	.av_readdata_pre_42(\cpu_jtag_debug_module_translator|av_readdata_pre[4]~q ),
	.av_readdata_pre_43(\led_pio_s1_translator|av_readdata_pre[4]~q ),
	.av_readdata_pre_44(\sys_clk_timer_s1_translator|av_readdata_pre[4]~q ),
	.src_data_4(src_data_4),
	.av_readdata_pre_201(\cpu_jtag_debug_module_translator|av_readdata_pre[20]~q ),
	.src_payload5(src_payload5),
	.av_readdata_pre_12(\cpu_jtag_debug_module_translator|av_readdata_pre[12]~q ),
	.av_readdata_pre_121(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[12]~q ),
	.av_readdata_pre_122(\sys_clk_timer_s1_translator|av_readdata_pre[12]~q ),
	.src_payload6(src_payload6),
	.av_readdata_pre_28(\cpu_jtag_debug_module_translator|av_readdata_pre[28]~q ),
	.src_payload7(src_payload7),
	.av_readdata_pre_61(\switches_pio_s1_translator|av_readdata_pre[6]~q ),
	.av_readdata_pre_62(\cpu_jtag_debug_module_translator|av_readdata_pre[6]~q ),
	.av_readdata_pre_63(\led_pio_s1_translator|av_readdata_pre[6]~q ),
	.av_readdata_pre_64(\sys_clk_timer_s1_translator|av_readdata_pre[6]~q ),
	.src_data_6(src_data_6),
	.av_readdata_pre_221(\cpu_jtag_debug_module_translator|av_readdata_pre[22]~q ),
	.src_payload8(src_payload8),
	.av_readdata_pre_14(\cpu_jtag_debug_module_translator|av_readdata_pre[14]~q ),
	.av_readdata_pre_141(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[14]~q ),
	.av_readdata_pre_142(\sys_clk_timer_s1_translator|av_readdata_pre[14]~q ),
	.src_payload9(src_payload9),
	.av_readdata_pre_301(\cpu_jtag_debug_module_translator|av_readdata_pre[30]~q ),
	.src_payload10(src_payload10),
	.av_readdata_pre_71(\switches_pio_s1_translator|av_readdata_pre[7]~q ),
	.av_readdata_pre_72(\cpu_jtag_debug_module_translator|av_readdata_pre[7]~q ),
	.av_readdata_pre_73(\led_pio_s1_translator|av_readdata_pre[7]~q ),
	.av_readdata_pre_74(\sys_clk_timer_s1_translator|av_readdata_pre[7]~q ),
	.src_data_7(src_data_7),
	.av_readdata_pre_23(\cpu_jtag_debug_module_translator|av_readdata_pre[23]~q ),
	.src_payload11(src_payload11),
	.av_readdata_pre_15(\cpu_jtag_debug_module_translator|av_readdata_pre[15]~q ),
	.av_readdata_pre_151(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[15]~q ),
	.av_readdata_pre_152(\sys_clk_timer_s1_translator|av_readdata_pre[15]~q ),
	.src_payload12(src_payload12),
	.av_readdata_pre_31(\cpu_jtag_debug_module_translator|av_readdata_pre[31]~q ),
	.src_payload13(src_payload13),
	.av_readdata_pre_11(\cpu_jtag_debug_module_translator|av_readdata_pre[11]~q ),
	.av_readdata_pre_111(\sys_clk_timer_s1_translator|av_readdata_pre[11]~q ),
	.src_payload14(src_payload14),
	.av_readdata_pre_27(\cpu_jtag_debug_module_translator|av_readdata_pre[27]~q ),
	.src_payload15(src_payload15),
	.av_readdata_pre_10(\cpu_jtag_debug_module_translator|av_readdata_pre[10]~q ),
	.av_readdata_pre_101(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[10]~q ),
	.av_readdata_pre_102(\sys_clk_timer_s1_translator|av_readdata_pre[10]~q ),
	.src_payload16(src_payload16),
	.av_readdata_pre_26(\cpu_jtag_debug_module_translator|av_readdata_pre[26]~q ),
	.src_payload17(src_payload17),
	.av_readdata_pre_25(\cpu_jtag_debug_module_translator|av_readdata_pre[25]~q ),
	.src_payload18(src_payload18),
	.av_readdata_pre_9(\led_pio_s1_translator|av_readdata_pre[9]~q ),
	.av_readdata_pre_91(\jtag_uart_avalon_jtag_slave_translator|av_readdata_pre[9]~q ),
	.av_readdata_pre_92(\sys_clk_timer_s1_translator|av_readdata_pre[9]~q ),
	.av_readdata_pre_93(\cpu_jtag_debug_module_translator|av_readdata_pre[9]~q ),
	.av_readdata_pre_94(\switches_pio_s1_translator|av_readdata_pre[9]~q ),
	.src_data_9(src_data_9),
	.av_readdata_pre_32(\led_pio_s1_translator|av_readdata_pre[3]~q ),
	.av_readdata_pre_33(\sys_clk_timer_s1_translator|av_readdata_pre[3]~q ),
	.av_readdata_pre_34(\cpu_jtag_debug_module_translator|av_readdata_pre[3]~q ),
	.av_readdata_pre_35(\switches_pio_s1_translator|av_readdata_pre[3]~q ),
	.src_data_3(src_data_3),
	.av_readdata_pre_191(\cpu_jtag_debug_module_translator|av_readdata_pre[19]~q ),
	.src_payload19(src_payload19),
	.av_readdata_pre_210(\led_pio_s1_translator|av_readdata_pre[2]~q ),
	.av_readdata_pre_212(\sys_clk_timer_s1_translator|av_readdata_pre[2]~q ),
	.av_readdata_pre_213(\cpu_jtag_debug_module_translator|av_readdata_pre[2]~q ),
	.av_readdata_pre_214(\switches_pio_s1_translator|av_readdata_pre[2]~q ),
	.src_data_2(src_data_2),
	.av_readdata_pre_181(\cpu_jtag_debug_module_translator|av_readdata_pre[18]~q ),
	.src_payload20(src_payload20),
	.av_readdata_pre_110(\led_pio_s1_translator|av_readdata_pre[1]~q ),
	.av_readdata_pre_112(\sys_clk_timer_s1_translator|av_readdata_pre[1]~q ),
	.av_readdata_pre_113(\cpu_jtag_debug_module_translator|av_readdata_pre[1]~q ),
	.av_readdata_pre_114(\switches_pio_s1_translator|av_readdata_pre[1]~q ),
	.src_data_1(src_data_1),
	.av_readdata_pre_171(\cpu_jtag_debug_module_translator|av_readdata_pre[17]~q ),
	.src_payload21(src_payload21));

processor_processor_mm_interconnect_0_rsp_demux_002_1 rsp_demux_003(
	.read_latency_shift_reg_0(\onchip_mem_s1_translator|read_latency_shift_reg[0]~q ),
	.mem_74_0(\onchip_mem_s1_agent_rsp_fifo|mem[0][74]~q ),
	.mem_56_0(\onchip_mem_s1_agent_rsp_fifo|mem[0][56]~q ),
	.src0_valid(\rsp_demux_003|src0_valid~0_combout ),
	.src1_valid(\rsp_demux_003|src1_valid~0_combout ));

processor_processor_mm_interconnect_0_rsp_demux_002 rsp_demux_002(
	.read_latency_shift_reg_0(\cpu_jtag_debug_module_translator|read_latency_shift_reg[0]~q ),
	.mem_74_0(\cpu_jtag_debug_module_agent_rsp_fifo|mem[0][74]~q ),
	.mem_56_0(\cpu_jtag_debug_module_agent_rsp_fifo|mem[0][56]~q ),
	.src0_valid(\rsp_demux_002|src0_valid~0_combout ),
	.src1_valid(\rsp_demux_002|src1_valid~0_combout ));

processor_processor_mm_interconnect_0_cmd_mux_002_1 cmd_mux_003(
	.M_st_data_8(M_st_data_8),
	.M_st_data_9(M_st_data_9),
	.M_st_data_16(M_st_data_16),
	.M_st_data_21(M_st_data_21),
	.M_st_data_13(M_st_data_13),
	.M_st_data_20(M_st_data_20),
	.M_st_data_12(M_st_data_12),
	.M_st_data_22(M_st_data_22),
	.M_st_data_14(M_st_data_14),
	.M_st_data_23(M_st_data_23),
	.M_st_data_15(M_st_data_15),
	.M_st_data_11(M_st_data_11),
	.M_st_data_10(M_st_data_10),
	.M_st_data_19(M_st_data_19),
	.M_st_data_18(M_st_data_18),
	.M_st_data_17(M_st_data_17),
	.M_st_data_0(M_st_data_0),
	.r_sync_rst(r_sync_rst),
	.M_alu_result_5(M_alu_result_5),
	.M_alu_result_4(M_alu_result_4),
	.M_alu_result_6(M_alu_result_6),
	.M_alu_result_14(M_alu_result_14),
	.M_alu_result_13(M_alu_result_13),
	.M_alu_result_12(M_alu_result_12),
	.M_alu_result_11(M_alu_result_11),
	.M_alu_result_10(M_alu_result_10),
	.M_alu_result_9(M_alu_result_9),
	.M_alu_result_8(M_alu_result_8),
	.M_alu_result_7(M_alu_result_7),
	.M_alu_result_3(M_alu_result_3),
	.M_alu_result_2(M_alu_result_2),
	.M_st_data_1(M_st_data_1),
	.M_st_data_2(M_st_data_2),
	.M_st_data_3(M_st_data_3),
	.M_st_data_4(M_st_data_4),
	.M_st_data_5(M_st_data_5),
	.M_st_data_6(M_st_data_6),
	.M_st_data_7(M_st_data_7),
	.saved_grant_0(saved_grant_01),
	.read_latency_shift_reg(\onchip_mem_s1_translator|read_latency_shift_reg~0_combout ),
	.ic_fill_tag_3(ic_fill_tag_3),
	.ic_fill_tag_2(ic_fill_tag_2),
	.ic_fill_tag_1(ic_fill_tag_1),
	.ic_fill_tag_0(ic_fill_tag_0),
	.src3_valid(src3_valid),
	.saved_grant_1(saved_grant_11),
	.src1_valid(src1_valid),
	.ic_fill_line_5(ic_fill_line_5),
	.ic_fill_line_0(ic_fill_line_0),
	.ic_fill_line_1(ic_fill_line_1),
	.ic_fill_line_2(ic_fill_line_2),
	.ic_fill_line_3(ic_fill_line_3),
	.ic_fill_line_4(ic_fill_line_4),
	.src_payload(src_payload22),
	.ic_fill_ap_offset_0(ic_fill_ap_offset_0),
	.src_data_38(src_data_38),
	.ic_fill_ap_offset_1(ic_fill_ap_offset_1),
	.src_data_39(src_data_39),
	.ic_fill_ap_offset_2(ic_fill_ap_offset_2),
	.src_data_40(src_data_40),
	.src_data_41(src_data_41),
	.src_data_42(src_data_42),
	.src_data_43(src_data_43),
	.src_data_44(src_data_44),
	.src_data_45(src_data_45),
	.src_data_46(src_data_461),
	.src_data_47(src_data_47),
	.src_data_48(src_data_48),
	.src_data_49(src_data_49),
	.src_data_50(src_data_50),
	.M_mem_byte_en_0(M_mem_byte_en_0),
	.src_data_32(src_data_32),
	.src_payload1(src_payload23),
	.M_mem_byte_en_2(M_mem_byte_en_2),
	.src_data_34(src_data_34),
	.src_payload2(src_payload24),
	.M_mem_byte_en_1(M_mem_byte_en_1),
	.src_data_33(src_data_33),
	.M_st_data_24(M_st_data_24),
	.src_payload3(src_payload25),
	.M_mem_byte_en_3(M_mem_byte_en_3),
	.src_data_35(src_data_35),
	.src_payload4(src_payload28),
	.src_payload5(src_payload29),
	.src_payload6(src_payload30),
	.M_st_data_29(M_st_data_29),
	.src_payload7(src_payload31),
	.src_payload8(src_payload32),
	.src_payload9(src_payload33),
	.src_payload10(src_payload34),
	.M_st_data_28(M_st_data_28),
	.src_payload11(src_payload35),
	.src_payload12(src_payload36),
	.src_payload13(src_payload37),
	.src_payload14(src_payload38),
	.M_st_data_30(M_st_data_30),
	.src_payload15(src_payload39),
	.src_payload16(src_payload40),
	.src_payload17(src_payload41),
	.src_payload18(src_payload42),
	.M_st_data_31(M_st_data_31),
	.src_payload19(src_payload43),
	.src_payload20(src_payload44),
	.M_st_data_27(M_st_data_27),
	.src_payload21(src_payload45),
	.src_payload22(src_payload46),
	.M_st_data_26(M_st_data_26),
	.src_payload23(src_payload47),
	.M_st_data_25(M_st_data_25),
	.src_payload24(src_payload48),
	.src_payload25(src_payload49),
	.src_payload26(src_payload50),
	.src_payload27(src_payload51),
	.src_payload28(src_payload52),
	.src_payload29(src_payload53),
	.src_payload30(src_payload54),
	.src_payload31(src_payload55),
	.clk_clk(clk_clk));

processor_processor_mm_interconnect_0_cmd_mux_002 cmd_mux_002(
	.M_st_data_8(M_st_data_8),
	.M_st_data_9(M_st_data_9),
	.M_st_data_16(M_st_data_16),
	.M_st_data_21(M_st_data_21),
	.M_st_data_13(M_st_data_13),
	.M_st_data_20(M_st_data_20),
	.M_st_data_12(M_st_data_12),
	.M_st_data_22(M_st_data_22),
	.M_st_data_14(M_st_data_14),
	.M_st_data_23(M_st_data_23),
	.M_st_data_15(M_st_data_15),
	.M_st_data_11(M_st_data_11),
	.M_st_data_10(M_st_data_10),
	.M_st_data_19(M_st_data_19),
	.M_st_data_18(M_st_data_18),
	.M_st_data_17(M_st_data_17),
	.M_st_data_0(M_st_data_0),
	.r_sync_rst(r_sync_rst),
	.M_alu_result_5(M_alu_result_5),
	.M_alu_result_4(M_alu_result_4),
	.M_alu_result_6(M_alu_result_6),
	.M_alu_result_10(M_alu_result_10),
	.M_alu_result_9(M_alu_result_9),
	.M_alu_result_8(M_alu_result_8),
	.M_alu_result_7(M_alu_result_7),
	.M_alu_result_3(M_alu_result_3),
	.M_alu_result_2(M_alu_result_2),
	.M_st_data_1(M_st_data_1),
	.M_st_data_2(M_st_data_2),
	.M_st_data_3(M_st_data_3),
	.M_st_data_4(M_st_data_4),
	.M_st_data_5(M_st_data_5),
	.M_st_data_6(M_st_data_6),
	.M_st_data_7(M_st_data_7),
	.saved_grant_0(saved_grant_0),
	.write(\cpu_jtag_debug_module_agent_rsp_fifo|write~0_combout ),
	.hbreak_enabled(hbreak_enabled),
	.src2_valid(src2_valid),
	.saved_grant_1(saved_grant_1),
	.src0_valid(src0_valid),
	.ic_fill_line_5(ic_fill_line_5),
	.src_data_46(src_data_46),
	.ic_fill_line_0(ic_fill_line_0),
	.ic_fill_line_1(ic_fill_line_1),
	.ic_fill_line_2(ic_fill_line_2),
	.ic_fill_line_3(ic_fill_line_3),
	.ic_fill_line_4(ic_fill_line_4),
	.ic_fill_ap_offset_0(ic_fill_ap_offset_0),
	.ic_fill_ap_offset_1(ic_fill_ap_offset_1),
	.ic_fill_ap_offset_2(ic_fill_ap_offset_2),
	.M_mem_byte_en_0(M_mem_byte_en_0),
	.M_mem_byte_en_2(M_mem_byte_en_2),
	.M_mem_byte_en_1(M_mem_byte_en_1),
	.M_st_data_24(M_st_data_24),
	.M_mem_byte_en_3(M_mem_byte_en_3),
	.src_payload(src_payload26),
	.src_data_38(src_data_381),
	.src_data_41(src_data_411),
	.src_data_40(src_data_401),
	.src_data_39(src_data_391),
	.src_data_45(src_data_451),
	.src_data_44(src_data_441),
	.src_data_43(src_data_431),
	.src_data_42(src_data_421),
	.src_payload1(src_payload27),
	.M_st_data_29(M_st_data_29),
	.M_st_data_28(M_st_data_28),
	.M_st_data_30(M_st_data_30),
	.M_st_data_31(M_st_data_31),
	.M_st_data_27(M_st_data_27),
	.M_st_data_26(M_st_data_26),
	.M_st_data_25(M_st_data_25),
	.src_payload2(src_payload56),
	.src_data_32(src_data_321),
	.src_payload3(src_payload57),
	.src_payload4(src_payload58),
	.src_payload5(src_payload59),
	.src_data_34(src_data_341),
	.src_payload6(src_payload60),
	.src_data_33(src_data_331),
	.src_payload7(src_payload61),
	.src_data_35(src_data_351),
	.src_payload8(src_payload62),
	.src_payload9(src_payload63),
	.src_payload10(src_payload64),
	.src_payload11(src_payload65),
	.src_payload12(src_payload66),
	.src_payload13(src_payload67),
	.src_payload14(src_payload68),
	.src_payload15(src_payload69),
	.src_payload16(src_payload70),
	.src_payload17(src_payload71),
	.src_payload18(src_payload72),
	.src_payload19(src_payload73),
	.src_payload20(src_payload74),
	.src_payload21(src_payload75),
	.src_payload22(src_payload76),
	.src_payload23(src_payload77),
	.src_payload24(src_payload78),
	.src_payload25(src_payload79),
	.src_payload26(src_payload80),
	.src_payload27(src_payload81),
	.src_payload28(src_payload82),
	.src_payload29(src_payload83),
	.src_payload30(src_payload84),
	.src_payload31(src_payload85),
	.src_payload32(src_payload86),
	.clk_clk(clk_clk));

processor_processor_mm_interconnect_0_cmd_demux_001 cmd_demux_001(
	.clr_break_line(clr_break_line),
	.write(\cpu_jtag_debug_module_agent_rsp_fifo|write~0_combout ),
	.read_latency_shift_reg(\onchip_mem_s1_translator|read_latency_shift_reg~0_combout ),
	.saved_grant_1(saved_grant_1),
	.i_read(i_read),
	.last_channel_0(\cpu_instruction_master_limiter|last_channel[0]~q ),
	.has_pending_responses(has_pending_responses),
	.Equal1(Equal11),
	.src0_valid(src0_valid),
	.saved_grant_11(saved_grant_11),
	.last_dest_id_1(last_dest_id_1),
	.src1_valid(src1_valid),
	.WideOr0(WideOr0));

processor_processor_mm_interconnect_0_cmd_demux cmd_demux(
	.clr_break_line(clr_break_line),
	.d_write(d_write),
	.Equal1(Equal1),
	.Equal2(Equal2),
	.Equal4(Equal4),
	.d_read(d_read),
	.mem_used_1(\sysid_control_slave_agent_rsp_fifo|mem_used[1]~q ),
	.read_accepted(read_accepted),
	.always1(\router|always1~0_combout ),
	.always11(\router|always1~1_combout ),
	.sink_ready(\cmd_demux|sink_ready~0_combout ),
	.wait_latency_counter_1(\sysid_control_slave_translator|wait_latency_counter[1]~q ),
	.wait_latency_counter_0(\sysid_control_slave_translator|wait_latency_counter[0]~q ),
	.sink_ready1(\cmd_demux|sink_ready~1_combout ),
	.mem_used_11(\switches_pio_s1_agent_rsp_fifo|mem_used[1]~q ),
	.always12(\router|always1~2_combout ),
	.sink_ready2(\cmd_demux|sink_ready~2_combout ),
	.wait_latency_counter_11(\switches_pio_s1_translator|wait_latency_counter[1]~q ),
	.wait_latency_counter_01(\switches_pio_s1_translator|wait_latency_counter[0]~q ),
	.sink_ready3(\cmd_demux|sink_ready~3_combout ),
	.Equal21(\router|Equal2~1_combout ),
	.mem_used_12(\jtag_uart_avalon_jtag_slave_agent_rsp_fifo|mem_used[1]~q ),
	.av_waitrequest(av_waitrequest),
	.Equal6(Equal6),
	.sink_ready4(\cmd_demux|sink_ready~4_combout ),
	.saved_grant_0(saved_grant_0),
	.write(\cpu_jtag_debug_module_agent_rsp_fifo|write~0_combout ),
	.saved_grant_01(saved_grant_01),
	.read_latency_shift_reg(\onchip_mem_s1_translator|read_latency_shift_reg~0_combout ),
	.Equal11(\router|Equal1~1_combout ),
	.WideOr0(\cmd_demux|WideOr0~0_combout ),
	.src2_valid(\cmd_demux|src2_valid~0_combout ),
	.src2_valid1(\cmd_demux|src2_valid~1_combout ),
	.src2_valid2(src2_valid),
	.src3_valid(src3_valid),
	.sink_ready5(\cmd_demux|sink_ready~5_combout ),
	.sink_ready6(\cmd_demux|sink_ready~6_combout ),
	.sink_ready7(\cmd_demux|sink_ready~7_combout ),
	.sink_ready8(\cmd_demux|sink_ready~8_combout ));

processor_altera_merlin_traffic_limiter cpu_instruction_master_limiter(
	.reset(r_sync_rst),
	.clr_break_line(clr_break_line),
	.i_read(i_read),
	.last_channel_0(\cpu_instruction_master_limiter|last_channel[0]~q ),
	.has_pending_responses1(has_pending_responses),
	.cmd_sink_channel({gnd,gnd,gnd,gnd,gnd,gnd,Equal11}),
	.last_dest_id_1(last_dest_id_1),
	.WideOr0(WideOr0),
	.nonposted_cmd_accepted1(nonposted_cmd_accepted),
	.src1_valid(\rsp_demux_002|src1_valid~0_combout ),
	.src1_valid1(\rsp_demux_003|src1_valid~0_combout ),
	.mem_61_0(\cpu_jtag_debug_module_agent_rsp_fifo|mem[0][61]~q ),
	.mem_61_01(\onchip_mem_s1_agent_rsp_fifo|mem[0][61]~q ),
	.clk(clk_clk));

processor_processor_mm_interconnect_0_router_001 router_001(
	.ic_fill_tag_5(ic_fill_tag_5),
	.ic_fill_tag_4(ic_fill_tag_4),
	.ic_fill_tag_3(ic_fill_tag_3),
	.ic_fill_tag_2(ic_fill_tag_2),
	.ic_fill_tag_1(ic_fill_tag_1),
	.ic_fill_tag_0(ic_fill_tag_0),
	.Equal1(Equal11));

processor_processor_mm_interconnect_0_router router(
	.M_alu_result_5(M_alu_result_5),
	.M_alu_result_4(M_alu_result_4),
	.M_alu_result_6(M_alu_result_6),
	.M_alu_result_16(M_alu_result_16),
	.M_alu_result_15(M_alu_result_15),
	.M_alu_result_14(M_alu_result_14),
	.M_alu_result_13(M_alu_result_13),
	.Equal1(Equal1),
	.M_alu_result_12(M_alu_result_12),
	.M_alu_result_11(M_alu_result_11),
	.M_alu_result_10(M_alu_result_10),
	.M_alu_result_9(M_alu_result_9),
	.M_alu_result_8(M_alu_result_8),
	.M_alu_result_7(M_alu_result_7),
	.Equal2(Equal2),
	.Equal4(Equal4),
	.M_alu_result_3(M_alu_result_3),
	.d_read(d_read),
	.read_accepted(read_accepted),
	.always1(\router|always1~0_combout ),
	.always11(\router|always1~1_combout ),
	.always12(\router|always1~2_combout ),
	.Equal21(\router|Equal2~1_combout ),
	.Equal6(Equal6),
	.Equal11(\router|Equal1~1_combout ),
	.Equal61(\router|Equal6~1_combout ));

processor_altera_avalon_sc_fifo_4 switches_pio_s1_agent_rsp_fifo(
	.reset(r_sync_rst),
	.read_latency_shift_reg_0(\switches_pio_s1_translator|read_latency_shift_reg[0]~q ),
	.mem_used_1(\switches_pio_s1_agent_rsp_fifo|mem_used[1]~q ),
	.sink_ready(\cmd_demux|sink_ready~3_combout ),
	.sink_ready1(\cmd_demux|sink_ready~7_combout ),
	.sink_ready2(\cmd_demux|sink_ready~8_combout ),
	.clk(clk_clk));

processor_altera_avalon_sc_fifo_2 led_pio_s1_agent_rsp_fifo(
	.reset(r_sync_rst),
	.clr_break_line(clr_break_line),
	.mem_used_1(mem_used_1),
	.Equal4(Equal4),
	.wait_latency_counter_1(wait_latency_counter_1),
	.read_latency_shift_reg_0(\led_pio_s1_translator|read_latency_shift_reg[0]~q ),
	.uav_read(uav_read),
	.av_waitrequest_generated(\led_pio_s1_translator|av_waitrequest_generated~0_combout ),
	.mem_used_11(\led_pio_s1_agent_rsp_fifo|mem_used[1]~0_combout ),
	.clk(clk_clk));

processor_altera_avalon_sc_fifo_5 sys_clk_timer_s1_agent_rsp_fifo(
	.reset(r_sync_rst),
	.clr_break_line(clr_break_line),
	.d_write(d_write),
	.read_latency_shift_reg_0(\sys_clk_timer_s1_translator|read_latency_shift_reg[0]~q ),
	.Equal2(\router|Equal2~1_combout ),
	.mem_used_1(mem_used_11),
	.wait_latency_counter_1(wait_latency_counter_11),
	.wait_latency_counter_0(wait_latency_counter_01),
	.uav_read(uav_read),
	.period_l_wr_strobe(period_l_wr_strobe),
	.mem_used_11(\sys_clk_timer_s1_agent_rsp_fifo|mem_used[1]~0_combout ),
	.read_latency_shift_reg(\sys_clk_timer_s1_translator|read_latency_shift_reg~0_combout ),
	.clk(clk_clk));

processor_altera_avalon_sc_fifo_3 onchip_mem_s1_agent_rsp_fifo(
	.reset(r_sync_rst),
	.clr_break_line(clr_break_line),
	.read_latency_shift_reg_0(\onchip_mem_s1_translator|read_latency_shift_reg[0]~q ),
	.mem_74_0(\onchip_mem_s1_agent_rsp_fifo|mem[0][74]~q ),
	.mem_56_0(\onchip_mem_s1_agent_rsp_fifo|mem[0][56]~q ),
	.saved_grant_0(saved_grant_01),
	.mem_used_1(mem_used_13),
	.uav_read(uav_read),
	.i_read(i_read),
	.saved_grant_1(saved_grant_11),
	.rf_source_valid(\onchip_mem_s1_agent|rf_source_valid~0_combout ),
	.read_latency_shift_reg(\onchip_mem_s1_translator|read_latency_shift_reg~1_combout ),
	.mem_61_0(\onchip_mem_s1_agent_rsp_fifo|mem[0][61]~q ),
	.clk(clk_clk));

endmodule

module processor_altera_avalon_sc_fifo (
	reset,
	read_latency_shift_reg_0,
	mem_74_0,
	mem_56_0,
	saved_grant_0,
	waitrequest,
	mem_used_1,
	write,
	uav_read,
	saved_grant_1,
	i_read,
	rf_source_valid,
	mem_61_0,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset;
input 	read_latency_shift_reg_0;
output 	mem_74_0;
output 	mem_56_0;
input 	saved_grant_0;
input 	waitrequest;
output 	mem_used_1;
output 	write;
input 	uav_read;
input 	saved_grant_1;
input 	i_read;
input 	rf_source_valid;
output 	mem_61_0;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \mem[1][74]~q ;
wire \mem~0_combout ;
wire \mem_used[0]~2_combout ;
wire \mem_used[0]~q ;
wire \mem_used[1]~0_combout ;
wire \mem[1][56]~q ;
wire \mem~1_combout ;
wire \mem_used[1]~1_combout ;
wire \mem[1][94]~q ;
wire \mem~2_combout ;


dffeas \mem[0][74] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[1]~0_combout ),
	.q(mem_74_0),
	.prn(vcc));
defparam \mem[0][74] .is_wysiwyg = "true";
defparam \mem[0][74] .power_up = "low";

dffeas \mem[0][56] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[1]~0_combout ),
	.q(mem_56_0),
	.prn(vcc));
defparam \mem[0][56] .is_wysiwyg = "true";
defparam \mem[0][56] .power_up = "low";

dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_1),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

cyclonev_lcell_comb \write~0 (
	.dataa(!waitrequest),
	.datab(!mem_used_1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(write),
	.sumout(),
	.cout(),
	.shareout());
defparam \write~0 .extended_lut = "off";
defparam \write~0 .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \write~0 .shared_arith = "off";

dffeas \mem[0][61] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[1]~0_combout ),
	.q(mem_61_0),
	.prn(vcc));
defparam \mem[0][61] .is_wysiwyg = "true";
defparam \mem[0][61] .power_up = "low";

dffeas \mem[1][74] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][74]~q ),
	.prn(vcc));
defparam \mem[1][74] .is_wysiwyg = "true";
defparam \mem[1][74] .power_up = "low";

cyclonev_lcell_comb \mem~0 (
	.dataa(!mem_used_1),
	.datab(!saved_grant_1),
	.datac(!\mem[1][74]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~0 .extended_lut = "off";
defparam \mem~0 .lut_mask = 64'h2727272727272727;
defparam \mem~0 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[0]~2 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!waitrequest),
	.datac(!mem_used_1),
	.datad(!rf_source_valid),
	.datae(!\mem_used[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[0]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[0]~2 .extended_lut = "off";
defparam \mem_used[0]~2 .lut_mask = 64'hACFFFFFFACFFFFFF;
defparam \mem_used[0]~2 .shared_arith = "off";

dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_used[0]~q ),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

cyclonev_lcell_comb \mem_used[1]~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!\mem_used[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~0 .extended_lut = "off";
defparam \mem_used[1]~0 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \mem_used[1]~0 .shared_arith = "off";

dffeas \mem[1][56] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][56]~q ),
	.prn(vcc));
defparam \mem[1][56] .is_wysiwyg = "true";
defparam \mem[1][56] .power_up = "low";

cyclonev_lcell_comb \mem~1 (
	.dataa(!uav_read),
	.datab(!saved_grant_0),
	.datac(!mem_used_1),
	.datad(!saved_grant_1),
	.datae(!i_read),
	.dataf(!\mem[1][56]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~1 .extended_lut = "off";
defparam \mem~1 .lut_mask = 64'h53FFFFFFFFFFFFFF;
defparam \mem~1 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[1]~1 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!waitrequest),
	.datac(!mem_used_1),
	.datad(!rf_source_valid),
	.datae(!\mem_used[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~1 .extended_lut = "off";
defparam \mem_used[1]~1 .lut_mask = 64'hAFFFCFFFAFFFCFFF;
defparam \mem_used[1]~1 .shared_arith = "off";

dffeas \mem[1][94] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][94]~q ),
	.prn(vcc));
defparam \mem[1][94] .is_wysiwyg = "true";
defparam \mem[1][94] .power_up = "low";

cyclonev_lcell_comb \mem~2 (
	.dataa(!saved_grant_0),
	.datab(!mem_used_1),
	.datac(!saved_grant_1),
	.datad(!\mem[1][94]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~2 .extended_lut = "off";
defparam \mem~2 .lut_mask = 64'h47FF47FF47FF47FF;
defparam \mem~2 .shared_arith = "off";

endmodule

module processor_altera_avalon_sc_fifo_1 (
	reset,
	clr_break_line,
	read_latency_shift_reg_0,
	mem_used_1,
	av_waitrequest,
	uav_read,
	Equal6,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset;
input 	clr_break_line;
input 	read_latency_shift_reg_0;
output 	mem_used_1;
input 	av_waitrequest;
input 	uav_read;
input 	Equal6;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \write~0_combout ;
wire \mem_used[0]~1_combout ;
wire \mem_used[0]~q ;
wire \mem_used[1]~0_combout ;


dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_1),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

cyclonev_lcell_comb \write~0 (
	.dataa(!clr_break_line),
	.datab(!av_waitrequest),
	.datac(!Equal6),
	.datad(!uav_read),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\write~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \write~0 .extended_lut = "off";
defparam \write~0 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \write~0 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[0]~1 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_1),
	.datac(!\mem_used[0]~q ),
	.datad(!\write~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[0]~1 .extended_lut = "off";
defparam \mem_used[0]~1 .lut_mask = 64'h8BFF8BFF8BFF8BFF;
defparam \mem_used[0]~1 .shared_arith = "off";

dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_used[0]~q ),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

cyclonev_lcell_comb \mem_used[1]~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_1),
	.datac(!\mem_used[0]~q ),
	.datad(!\write~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~0 .extended_lut = "off";
defparam \mem_used[1]~0 .lut_mask = 64'hA3FFA3FFA3FFA3FF;
defparam \mem_used[1]~0 .shared_arith = "off";

endmodule

module processor_altera_avalon_sc_fifo_2 (
	reset,
	clr_break_line,
	mem_used_1,
	Equal4,
	wait_latency_counter_1,
	read_latency_shift_reg_0,
	uav_read,
	av_waitrequest_generated,
	mem_used_11,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset;
input 	clr_break_line;
output 	mem_used_1;
input 	Equal4;
input 	wait_latency_counter_1;
input 	read_latency_shift_reg_0;
input 	uav_read;
input 	av_waitrequest_generated;
output 	mem_used_11;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \mem_used[0]~2_combout ;
wire \mem_used[0]~q ;
wire \mem_used[1]~1_combout ;


dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_1),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

cyclonev_lcell_comb \mem_used[1]~0 (
	.dataa(!wait_latency_counter_1),
	.datab(!clr_break_line),
	.datac(!Equal4),
	.datad(!uav_read),
	.datae(!av_waitrequest_generated),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(mem_used_11),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~0 .extended_lut = "off";
defparam \mem_used[1]~0 .lut_mask = 64'hBFFFFFFFBFFFFFFF;
defparam \mem_used[1]~0 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[0]~2 (
	.dataa(!mem_used_1),
	.datab(!read_latency_shift_reg_0),
	.datac(!\mem_used[0]~q ),
	.datad(!mem_used_11),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[0]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[0]~2 .extended_lut = "off";
defparam \mem_used[0]~2 .lut_mask = 64'h8DFF8DFF8DFF8DFF;
defparam \mem_used[0]~2 .shared_arith = "off";

dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_used[0]~q ),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

cyclonev_lcell_comb \mem_used[1]~1 (
	.dataa(!mem_used_1),
	.datab(!read_latency_shift_reg_0),
	.datac(!\mem_used[0]~q ),
	.datad(!mem_used_11),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~1 .extended_lut = "off";
defparam \mem_used[1]~1 .lut_mask = 64'hC5FFC5FFC5FFC5FF;
defparam \mem_used[1]~1 .shared_arith = "off";

endmodule

module processor_altera_avalon_sc_fifo_3 (
	reset,
	clr_break_line,
	read_latency_shift_reg_0,
	mem_74_0,
	mem_56_0,
	saved_grant_0,
	mem_used_1,
	uav_read,
	i_read,
	saved_grant_1,
	rf_source_valid,
	read_latency_shift_reg,
	mem_61_0,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset;
input 	clr_break_line;
input 	read_latency_shift_reg_0;
output 	mem_74_0;
output 	mem_56_0;
input 	saved_grant_0;
output 	mem_used_1;
input 	uav_read;
input 	i_read;
input 	saved_grant_1;
input 	rf_source_valid;
input 	read_latency_shift_reg;
output 	mem_61_0;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \mem[1][74]~q ;
wire \mem~0_combout ;
wire \mem_used[0]~2_combout ;
wire \mem_used[0]~q ;
wire \mem_used[1]~0_combout ;
wire \mem[1][56]~q ;
wire \mem~1_combout ;
wire \mem_used[1]~1_combout ;
wire \mem[1][94]~q ;
wire \mem~2_combout ;


dffeas \mem[0][74] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[1]~0_combout ),
	.q(mem_74_0),
	.prn(vcc));
defparam \mem[0][74] .is_wysiwyg = "true";
defparam \mem[0][74] .power_up = "low";

dffeas \mem[0][56] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[1]~0_combout ),
	.q(mem_56_0),
	.prn(vcc));
defparam \mem[0][56] .is_wysiwyg = "true";
defparam \mem[0][56] .power_up = "low";

dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_1),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

dffeas \mem[0][61] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[1]~0_combout ),
	.q(mem_61_0),
	.prn(vcc));
defparam \mem[0][61] .is_wysiwyg = "true";
defparam \mem[0][61] .power_up = "low";

dffeas \mem[1][74] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][74]~q ),
	.prn(vcc));
defparam \mem[1][74] .is_wysiwyg = "true";
defparam \mem[1][74] .power_up = "low";

cyclonev_lcell_comb \mem~0 (
	.dataa(!mem_used_1),
	.datab(!saved_grant_1),
	.datac(!\mem[1][74]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~0 .extended_lut = "off";
defparam \mem~0 .lut_mask = 64'h2727272727272727;
defparam \mem~0 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[0]~2 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_1),
	.datac(!read_latency_shift_reg),
	.datad(!\mem_used[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[0]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[0]~2 .extended_lut = "off";
defparam \mem_used[0]~2 .lut_mask = 64'hBFFFBFFFBFFFBFFF;
defparam \mem_used[0]~2 .shared_arith = "off";

dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_used[0]~q ),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

cyclonev_lcell_comb \mem_used[1]~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!\mem_used[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~0 .extended_lut = "off";
defparam \mem_used[1]~0 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \mem_used[1]~0 .shared_arith = "off";

dffeas \mem[1][56] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][56]~q ),
	.prn(vcc));
defparam \mem[1][56] .is_wysiwyg = "true";
defparam \mem[1][56] .power_up = "low";

cyclonev_lcell_comb \mem~1 (
	.dataa(!uav_read),
	.datab(!saved_grant_0),
	.datac(!mem_used_1),
	.datad(!i_read),
	.datae(!saved_grant_1),
	.dataf(!\mem[1][56]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~1 .extended_lut = "off";
defparam \mem~1 .lut_mask = 64'h53FFFFFFFFFFFFFF;
defparam \mem~1 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[1]~1 (
	.dataa(!clr_break_line),
	.datab(!read_latency_shift_reg_0),
	.datac(!mem_used_1),
	.datad(!rf_source_valid),
	.datae(!\mem_used[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~1 .extended_lut = "off";
defparam \mem_used[1]~1 .lut_mask = 64'hCFFF5FFFCFFF5FFF;
defparam \mem_used[1]~1 .shared_arith = "off";

dffeas \mem[1][94] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][94]~q ),
	.prn(vcc));
defparam \mem[1][94] .is_wysiwyg = "true";
defparam \mem[1][94] .power_up = "low";

cyclonev_lcell_comb \mem~2 (
	.dataa(!saved_grant_0),
	.datab(!mem_used_1),
	.datac(!saved_grant_1),
	.datad(!\mem[1][94]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~2 .extended_lut = "off";
defparam \mem~2 .lut_mask = 64'h47FF47FF47FF47FF;
defparam \mem~2 .shared_arith = "off";

endmodule

module processor_altera_avalon_sc_fifo_4 (
	reset,
	read_latency_shift_reg_0,
	mem_used_1,
	sink_ready,
	sink_ready1,
	sink_ready2,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset;
input 	read_latency_shift_reg_0;
output 	mem_used_1;
input 	sink_ready;
input 	sink_ready1;
input 	sink_ready2;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \mem_used[0]~1_combout ;
wire \mem_used[0]~q ;
wire \mem_used[1]~0_combout ;


dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_1),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

cyclonev_lcell_comb \mem_used[0]~1 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_1),
	.datac(!sink_ready),
	.datad(!\mem_used[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[0]~1 .extended_lut = "off";
defparam \mem_used[0]~1 .lut_mask = 64'hBFFFBFFFBFFFBFFF;
defparam \mem_used[0]~1 .shared_arith = "off";

dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_used[0]~q ),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

cyclonev_lcell_comb \mem_used[1]~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_1),
	.datac(!sink_ready1),
	.datad(!sink_ready2),
	.datae(!\mem_used[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~0 .extended_lut = "off";
defparam \mem_used[1]~0 .lut_mask = 64'hAFFF3FFFAFFF3FFF;
defparam \mem_used[1]~0 .shared_arith = "off";

endmodule

module processor_altera_avalon_sc_fifo_5 (
	reset,
	clr_break_line,
	d_write,
	read_latency_shift_reg_0,
	Equal2,
	mem_used_1,
	wait_latency_counter_1,
	wait_latency_counter_0,
	uav_read,
	period_l_wr_strobe,
	mem_used_11,
	read_latency_shift_reg,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset;
input 	clr_break_line;
input 	d_write;
input 	read_latency_shift_reg_0;
input 	Equal2;
output 	mem_used_1;
input 	wait_latency_counter_1;
input 	wait_latency_counter_0;
input 	uav_read;
input 	period_l_wr_strobe;
output 	mem_used_11;
input 	read_latency_shift_reg;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \mem_used[0]~2_combout ;
wire \mem_used[0]~q ;
wire \mem_used[1]~1_combout ;


dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_1),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

cyclonev_lcell_comb \mem_used[1]~0 (
	.dataa(!d_write),
	.datab(!uav_read),
	.datac(!wait_latency_counter_1),
	.datad(!wait_latency_counter_0),
	.datae(!period_l_wr_strobe),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(mem_used_11),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~0 .extended_lut = "off";
defparam \mem_used[1]~0 .lut_mask = 64'hFBF7F7FBFBF7F7FB;
defparam \mem_used[1]~0 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[0]~2 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_1),
	.datac(!read_latency_shift_reg),
	.datad(!\mem_used[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[0]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[0]~2 .extended_lut = "off";
defparam \mem_used[0]~2 .lut_mask = 64'hBFFFBFFFBFFFBFFF;
defparam \mem_used[0]~2 .shared_arith = "off";

dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_used[0]~q ),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

cyclonev_lcell_comb \mem_used[1]~1 (
	.dataa(!clr_break_line),
	.datab(!read_latency_shift_reg_0),
	.datac(!Equal2),
	.datad(!mem_used_1),
	.datae(!mem_used_11),
	.dataf(!\mem_used[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~1 .extended_lut = "off";
defparam \mem_used[1]~1 .lut_mask = 64'hCFFFFFFF5FFFFFFF;
defparam \mem_used[1]~1 .shared_arith = "off";

endmodule

module processor_altera_avalon_sc_fifo_6 (
	reset,
	read_latency_shift_reg_0,
	mem_used_1,
	sink_ready,
	sink_ready1,
	sink_ready2,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset;
input 	read_latency_shift_reg_0;
output 	mem_used_1;
input 	sink_ready;
input 	sink_ready1;
input 	sink_ready2;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \mem_used[0]~1_combout ;
wire \mem_used[0]~q ;
wire \mem_used[1]~0_combout ;


dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_1),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

cyclonev_lcell_comb \mem_used[0]~1 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_1),
	.datac(!sink_ready),
	.datad(!\mem_used[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[0]~1 .extended_lut = "off";
defparam \mem_used[0]~1 .lut_mask = 64'hBFFFBFFFBFFFBFFF;
defparam \mem_used[0]~1 .shared_arith = "off";

dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_used[0]~q ),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

cyclonev_lcell_comb \mem_used[1]~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_used_1),
	.datac(!sink_ready1),
	.datad(!sink_ready2),
	.datae(!\mem_used[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~0 .extended_lut = "off";
defparam \mem_used[1]~0 .lut_mask = 64'hAFFF3FFFAFFF3FFF;
defparam \mem_used[1]~0 .shared_arith = "off";

endmodule

module processor_altera_merlin_master_translator (
	reset,
	clr_break_line,
	d_write,
	mem_used_1,
	Equal4,
	wait_latency_counter_1,
	wait_latency_counter_0,
	d_read,
	WideOr1,
	read_accepted1,
	sink_ready,
	sink_ready1,
	Equal2,
	mem_used_11,
	wait_latency_counter_11,
	wait_latency_counter_01,
	sink_ready2,
	WideOr0,
	src2_valid,
	read_accepted2,
	uav_read,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset;
input 	clr_break_line;
input 	d_write;
input 	mem_used_1;
input 	Equal4;
input 	wait_latency_counter_1;
input 	wait_latency_counter_0;
input 	d_read;
input 	WideOr1;
output 	read_accepted1;
input 	sink_ready;
input 	sink_ready1;
input 	Equal2;
input 	mem_used_11;
input 	wait_latency_counter_11;
input 	wait_latency_counter_01;
input 	sink_ready2;
input 	WideOr0;
input 	src2_valid;
output 	read_accepted2;
output 	uav_read;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \read_accepted~1_combout ;
wire \read_accepted~2_combout ;
wire \read_accepted~3_combout ;
wire \read_accepted~4_combout ;
wire \read_accepted~5_combout ;


dffeas read_accepted(
	.clk(clk),
	.d(\read_accepted~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_accepted1),
	.prn(vcc));
defparam read_accepted.is_wysiwyg = "true";
defparam read_accepted.power_up = "low";

cyclonev_lcell_comb \read_accepted~0 (
	.dataa(!clr_break_line),
	.datab(!sink_ready),
	.datac(!sink_ready1),
	.datad(!sink_ready2),
	.datae(!\read_accepted~4_combout ),
	.dataf(!\read_accepted~5_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(read_accepted2),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_accepted~0 .extended_lut = "off";
defparam \read_accepted~0 .lut_mask = 64'hFFFFFFFFFFFF7FFF;
defparam \read_accepted~0 .shared_arith = "off";

cyclonev_lcell_comb \uav_read~0 (
	.dataa(!d_read),
	.datab(!read_accepted1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(uav_read),
	.sumout(),
	.cout(),
	.shareout());
defparam \uav_read~0 .extended_lut = "off";
defparam \uav_read~0 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \uav_read~0 .shared_arith = "off";

cyclonev_lcell_comb \read_accepted~1 (
	.dataa(!d_read),
	.datab(!WideOr1),
	.datac(!read_accepted1),
	.datad(!read_accepted2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_accepted~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_accepted~1 .extended_lut = "off";
defparam \read_accepted~1 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \read_accepted~1 .shared_arith = "off";

cyclonev_lcell_comb \read_accepted~2 (
	.dataa(!d_write),
	.datab(!mem_used_11),
	.datac(!wait_latency_counter_11),
	.datad(!wait_latency_counter_01),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_accepted~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_accepted~2 .extended_lut = "off";
defparam \read_accepted~2 .lut_mask = 64'hFDFEFDFEFDFEFDFE;
defparam \read_accepted~2 .shared_arith = "off";

cyclonev_lcell_comb \read_accepted~3 (
	.dataa(!wait_latency_counter_1),
	.datab(!wait_latency_counter_0),
	.datac(!d_write),
	.datad(!mem_used_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_accepted~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_accepted~3 .extended_lut = "off";
defparam \read_accepted~3 .lut_mask = 64'hFFBEFFBEFFBEFFBE;
defparam \read_accepted~3 .shared_arith = "off";

cyclonev_lcell_comb \read_accepted~4 (
	.dataa(!Equal4),
	.datab(!Equal2),
	.datac(!src2_valid),
	.datad(!\read_accepted~2_combout ),
	.datae(!\read_accepted~3_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_accepted~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_accepted~4 .extended_lut = "off";
defparam \read_accepted~4 .lut_mask = 64'hFFFFFF6FFFFFFF6F;
defparam \read_accepted~4 .shared_arith = "off";

cyclonev_lcell_comb \read_accepted~5 (
	.dataa(!Equal4),
	.datab(!WideOr0),
	.datac(!Equal2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_accepted~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_accepted~5 .extended_lut = "off";
defparam \read_accepted~5 .lut_mask = 64'hFEFEFEFEFEFEFEFE;
defparam \read_accepted~5 .shared_arith = "off";

endmodule

module processor_altera_merlin_slave_agent (
	saved_grant_0,
	uav_read,
	src2_valid,
	saved_grant_1,
	i_read,
	src0_valid,
	rf_source_valid)/* synthesis synthesis_greybox=1 */;
input 	saved_grant_0;
input 	uav_read;
input 	src2_valid;
input 	saved_grant_1;
input 	i_read;
input 	src0_valid;
output 	rf_source_valid;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb \rf_source_valid~0 (
	.dataa(!uav_read),
	.datab(!saved_grant_0),
	.datac(!src2_valid),
	.datad(!saved_grant_1),
	.datae(!i_read),
	.dataf(!src0_valid),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(rf_source_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \rf_source_valid~0 .extended_lut = "off";
defparam \rf_source_valid~0 .lut_mask = 64'h7FFFFFFFFFFFFFFF;
defparam \rf_source_valid~0 .shared_arith = "off";

endmodule

module processor_altera_merlin_slave_agent_3 (
	saved_grant_0,
	uav_read,
	i_read,
	src3_valid,
	saved_grant_1,
	src1_valid,
	rf_source_valid)/* synthesis synthesis_greybox=1 */;
input 	saved_grant_0;
input 	uav_read;
input 	i_read;
input 	src3_valid;
input 	saved_grant_1;
input 	src1_valid;
output 	rf_source_valid;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb \rf_source_valid~0 (
	.dataa(!uav_read),
	.datab(!saved_grant_0),
	.datac(!i_read),
	.datad(!src3_valid),
	.datae(!saved_grant_1),
	.dataf(!src1_valid),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(rf_source_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \rf_source_valid~0 .extended_lut = "off";
defparam \rf_source_valid~0 .lut_mask = 64'h7FFFFFFFFFFFFFFF;
defparam \rf_source_valid~0 .shared_arith = "off";

endmodule

module processor_altera_merlin_slave_translator (
	av_readdata,
	reset,
	clr_break_line,
	read_latency_shift_reg_0,
	write,
	rf_source_valid,
	av_readdata_pre_0,
	av_readdata_pre_16,
	av_readdata_pre_8,
	av_readdata_pre_24,
	av_readdata_pre_5,
	av_readdata_pre_21,
	av_readdata_pre_13,
	av_readdata_pre_29,
	av_readdata_pre_4,
	av_readdata_pre_20,
	av_readdata_pre_12,
	av_readdata_pre_28,
	av_readdata_pre_6,
	av_readdata_pre_22,
	av_readdata_pre_14,
	av_readdata_pre_30,
	av_readdata_pre_7,
	av_readdata_pre_23,
	av_readdata_pre_15,
	av_readdata_pre_31,
	av_readdata_pre_11,
	av_readdata_pre_27,
	av_readdata_pre_10,
	av_readdata_pre_26,
	av_readdata_pre_25,
	av_readdata_pre_9,
	av_readdata_pre_3,
	av_readdata_pre_19,
	av_readdata_pre_2,
	av_readdata_pre_18,
	av_readdata_pre_1,
	av_readdata_pre_17,
	clk)/* synthesis synthesis_greybox=1 */;
input 	[31:0] av_readdata;
input 	reset;
input 	clr_break_line;
output 	read_latency_shift_reg_0;
input 	write;
input 	rf_source_valid;
output 	av_readdata_pre_0;
output 	av_readdata_pre_16;
output 	av_readdata_pre_8;
output 	av_readdata_pre_24;
output 	av_readdata_pre_5;
output 	av_readdata_pre_21;
output 	av_readdata_pre_13;
output 	av_readdata_pre_29;
output 	av_readdata_pre_4;
output 	av_readdata_pre_20;
output 	av_readdata_pre_12;
output 	av_readdata_pre_28;
output 	av_readdata_pre_6;
output 	av_readdata_pre_22;
output 	av_readdata_pre_14;
output 	av_readdata_pre_30;
output 	av_readdata_pre_7;
output 	av_readdata_pre_23;
output 	av_readdata_pre_15;
output 	av_readdata_pre_31;
output 	av_readdata_pre_11;
output 	av_readdata_pre_27;
output 	av_readdata_pre_10;
output 	av_readdata_pre_26;
output 	av_readdata_pre_25;
output 	av_readdata_pre_9;
output 	av_readdata_pre_3;
output 	av_readdata_pre_19;
output 	av_readdata_pre_2;
output 	av_readdata_pre_18;
output 	av_readdata_pre_1;
output 	av_readdata_pre_17;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \read_latency_shift_reg~0_combout ;


dffeas \read_latency_shift_reg[0] (
	.clk(clk),
	.d(\read_latency_shift_reg~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_latency_shift_reg_0),
	.prn(vcc));
defparam \read_latency_shift_reg[0] .is_wysiwyg = "true";
defparam \read_latency_shift_reg[0] .power_up = "low";

dffeas \av_readdata_pre[0] (
	.clk(clk),
	.d(av_readdata[0]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_0),
	.prn(vcc));
defparam \av_readdata_pre[0] .is_wysiwyg = "true";
defparam \av_readdata_pre[0] .power_up = "low";

dffeas \av_readdata_pre[16] (
	.clk(clk),
	.d(av_readdata[16]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_16),
	.prn(vcc));
defparam \av_readdata_pre[16] .is_wysiwyg = "true";
defparam \av_readdata_pre[16] .power_up = "low";

dffeas \av_readdata_pre[8] (
	.clk(clk),
	.d(av_readdata[8]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_8),
	.prn(vcc));
defparam \av_readdata_pre[8] .is_wysiwyg = "true";
defparam \av_readdata_pre[8] .power_up = "low";

dffeas \av_readdata_pre[24] (
	.clk(clk),
	.d(av_readdata[24]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_24),
	.prn(vcc));
defparam \av_readdata_pre[24] .is_wysiwyg = "true";
defparam \av_readdata_pre[24] .power_up = "low";

dffeas \av_readdata_pre[5] (
	.clk(clk),
	.d(av_readdata[5]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_5),
	.prn(vcc));
defparam \av_readdata_pre[5] .is_wysiwyg = "true";
defparam \av_readdata_pre[5] .power_up = "low";

dffeas \av_readdata_pre[21] (
	.clk(clk),
	.d(av_readdata[21]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_21),
	.prn(vcc));
defparam \av_readdata_pre[21] .is_wysiwyg = "true";
defparam \av_readdata_pre[21] .power_up = "low";

dffeas \av_readdata_pre[13] (
	.clk(clk),
	.d(av_readdata[13]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_13),
	.prn(vcc));
defparam \av_readdata_pre[13] .is_wysiwyg = "true";
defparam \av_readdata_pre[13] .power_up = "low";

dffeas \av_readdata_pre[29] (
	.clk(clk),
	.d(av_readdata[29]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_29),
	.prn(vcc));
defparam \av_readdata_pre[29] .is_wysiwyg = "true";
defparam \av_readdata_pre[29] .power_up = "low";

dffeas \av_readdata_pre[4] (
	.clk(clk),
	.d(av_readdata[4]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_4),
	.prn(vcc));
defparam \av_readdata_pre[4] .is_wysiwyg = "true";
defparam \av_readdata_pre[4] .power_up = "low";

dffeas \av_readdata_pre[20] (
	.clk(clk),
	.d(av_readdata[20]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_20),
	.prn(vcc));
defparam \av_readdata_pre[20] .is_wysiwyg = "true";
defparam \av_readdata_pre[20] .power_up = "low";

dffeas \av_readdata_pre[12] (
	.clk(clk),
	.d(av_readdata[12]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_12),
	.prn(vcc));
defparam \av_readdata_pre[12] .is_wysiwyg = "true";
defparam \av_readdata_pre[12] .power_up = "low";

dffeas \av_readdata_pre[28] (
	.clk(clk),
	.d(av_readdata[28]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_28),
	.prn(vcc));
defparam \av_readdata_pre[28] .is_wysiwyg = "true";
defparam \av_readdata_pre[28] .power_up = "low";

dffeas \av_readdata_pre[6] (
	.clk(clk),
	.d(av_readdata[6]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_6),
	.prn(vcc));
defparam \av_readdata_pre[6] .is_wysiwyg = "true";
defparam \av_readdata_pre[6] .power_up = "low";

dffeas \av_readdata_pre[22] (
	.clk(clk),
	.d(av_readdata[22]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_22),
	.prn(vcc));
defparam \av_readdata_pre[22] .is_wysiwyg = "true";
defparam \av_readdata_pre[22] .power_up = "low";

dffeas \av_readdata_pre[14] (
	.clk(clk),
	.d(av_readdata[14]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_14),
	.prn(vcc));
defparam \av_readdata_pre[14] .is_wysiwyg = "true";
defparam \av_readdata_pre[14] .power_up = "low";

dffeas \av_readdata_pre[30] (
	.clk(clk),
	.d(av_readdata[30]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_30),
	.prn(vcc));
defparam \av_readdata_pre[30] .is_wysiwyg = "true";
defparam \av_readdata_pre[30] .power_up = "low";

dffeas \av_readdata_pre[7] (
	.clk(clk),
	.d(av_readdata[7]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_7),
	.prn(vcc));
defparam \av_readdata_pre[7] .is_wysiwyg = "true";
defparam \av_readdata_pre[7] .power_up = "low";

dffeas \av_readdata_pre[23] (
	.clk(clk),
	.d(av_readdata[23]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_23),
	.prn(vcc));
defparam \av_readdata_pre[23] .is_wysiwyg = "true";
defparam \av_readdata_pre[23] .power_up = "low";

dffeas \av_readdata_pre[15] (
	.clk(clk),
	.d(av_readdata[15]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_15),
	.prn(vcc));
defparam \av_readdata_pre[15] .is_wysiwyg = "true";
defparam \av_readdata_pre[15] .power_up = "low";

dffeas \av_readdata_pre[31] (
	.clk(clk),
	.d(av_readdata[31]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_31),
	.prn(vcc));
defparam \av_readdata_pre[31] .is_wysiwyg = "true";
defparam \av_readdata_pre[31] .power_up = "low";

dffeas \av_readdata_pre[11] (
	.clk(clk),
	.d(av_readdata[11]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_11),
	.prn(vcc));
defparam \av_readdata_pre[11] .is_wysiwyg = "true";
defparam \av_readdata_pre[11] .power_up = "low";

dffeas \av_readdata_pre[27] (
	.clk(clk),
	.d(av_readdata[27]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_27),
	.prn(vcc));
defparam \av_readdata_pre[27] .is_wysiwyg = "true";
defparam \av_readdata_pre[27] .power_up = "low";

dffeas \av_readdata_pre[10] (
	.clk(clk),
	.d(av_readdata[10]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_10),
	.prn(vcc));
defparam \av_readdata_pre[10] .is_wysiwyg = "true";
defparam \av_readdata_pre[10] .power_up = "low";

dffeas \av_readdata_pre[26] (
	.clk(clk),
	.d(av_readdata[26]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_26),
	.prn(vcc));
defparam \av_readdata_pre[26] .is_wysiwyg = "true";
defparam \av_readdata_pre[26] .power_up = "low";

dffeas \av_readdata_pre[25] (
	.clk(clk),
	.d(av_readdata[25]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_25),
	.prn(vcc));
defparam \av_readdata_pre[25] .is_wysiwyg = "true";
defparam \av_readdata_pre[25] .power_up = "low";

dffeas \av_readdata_pre[9] (
	.clk(clk),
	.d(av_readdata[9]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_9),
	.prn(vcc));
defparam \av_readdata_pre[9] .is_wysiwyg = "true";
defparam \av_readdata_pre[9] .power_up = "low";

dffeas \av_readdata_pre[3] (
	.clk(clk),
	.d(av_readdata[3]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_3),
	.prn(vcc));
defparam \av_readdata_pre[3] .is_wysiwyg = "true";
defparam \av_readdata_pre[3] .power_up = "low";

dffeas \av_readdata_pre[19] (
	.clk(clk),
	.d(av_readdata[19]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_19),
	.prn(vcc));
defparam \av_readdata_pre[19] .is_wysiwyg = "true";
defparam \av_readdata_pre[19] .power_up = "low";

dffeas \av_readdata_pre[2] (
	.clk(clk),
	.d(av_readdata[2]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_2),
	.prn(vcc));
defparam \av_readdata_pre[2] .is_wysiwyg = "true";
defparam \av_readdata_pre[2] .power_up = "low";

dffeas \av_readdata_pre[18] (
	.clk(clk),
	.d(av_readdata[18]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_18),
	.prn(vcc));
defparam \av_readdata_pre[18] .is_wysiwyg = "true";
defparam \av_readdata_pre[18] .power_up = "low";

dffeas \av_readdata_pre[1] (
	.clk(clk),
	.d(av_readdata[1]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_1),
	.prn(vcc));
defparam \av_readdata_pre[1] .is_wysiwyg = "true";
defparam \av_readdata_pre[1] .power_up = "low";

dffeas \av_readdata_pre[17] (
	.clk(clk),
	.d(av_readdata[17]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_17),
	.prn(vcc));
defparam \av_readdata_pre[17] .is_wysiwyg = "true";
defparam \av_readdata_pre[17] .power_up = "low";

cyclonev_lcell_comb \read_latency_shift_reg~0 (
	.dataa(!clr_break_line),
	.datab(!write),
	.datac(!rf_source_valid),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_latency_shift_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_latency_shift_reg~0 .extended_lut = "off";
defparam \read_latency_shift_reg~0 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \read_latency_shift_reg~0 .shared_arith = "off";

endmodule

module processor_altera_merlin_slave_translator_1 (
	av_readdata_pre_0,
	av_readdata_pre_16,
	av_readdata_pre_5,
	av_readdata_pre_21,
	av_readdata_pre_4,
	av_readdata_pre_20,
	av_readdata_pre_6,
	av_readdata_pre_22,
	av_readdata_pre_7,
	av_readdata_pre_3,
	av_readdata_pre_19,
	av_readdata_pre_2,
	av_readdata_pre_18,
	av_readdata_pre_1,
	av_readdata_pre_17,
	q_b_0,
	av_readdata,
	q_b_5,
	q_b_4,
	q_b_6,
	q_b_7,
	q_b_3,
	q_b_2,
	q_b_1,
	reset,
	clr_break_line,
	read_latency_shift_reg_0,
	mem_used_1,
	av_waitrequest,
	uav_read,
	Equal6,
	read_latency_shift_reg,
	av_readdata_pre_8,
	av_readdata_pre_13,
	av_readdata_pre_12,
	av_readdata_pre_14,
	av_readdata_pre_15,
	av_readdata_pre_10,
	av_readdata_pre_9,
	b_full,
	read_0,
	counter_reg_bit_0,
	counter_reg_bit_5,
	b_full1,
	counter_reg_bit_4,
	counter_reg_bit_3,
	counter_reg_bit_2,
	counter_reg_bit_1,
	clk)/* synthesis synthesis_greybox=1 */;
output 	av_readdata_pre_0;
output 	av_readdata_pre_16;
output 	av_readdata_pre_5;
output 	av_readdata_pre_21;
output 	av_readdata_pre_4;
output 	av_readdata_pre_20;
output 	av_readdata_pre_6;
output 	av_readdata_pre_22;
output 	av_readdata_pre_7;
output 	av_readdata_pre_3;
output 	av_readdata_pre_19;
output 	av_readdata_pre_2;
output 	av_readdata_pre_18;
output 	av_readdata_pre_1;
output 	av_readdata_pre_17;
input 	q_b_0;
input 	[31:0] av_readdata;
input 	q_b_5;
input 	q_b_4;
input 	q_b_6;
input 	q_b_7;
input 	q_b_3;
input 	q_b_2;
input 	q_b_1;
input 	reset;
input 	clr_break_line;
output 	read_latency_shift_reg_0;
input 	mem_used_1;
input 	av_waitrequest;
input 	uav_read;
input 	Equal6;
output 	read_latency_shift_reg;
output 	av_readdata_pre_8;
output 	av_readdata_pre_13;
output 	av_readdata_pre_12;
output 	av_readdata_pre_14;
output 	av_readdata_pre_15;
output 	av_readdata_pre_10;
output 	av_readdata_pre_9;
input 	b_full;
input 	read_0;
input 	counter_reg_bit_0;
input 	counter_reg_bit_5;
input 	b_full1;
input 	counter_reg_bit_4;
input 	counter_reg_bit_3;
input 	counter_reg_bit_2;
input 	counter_reg_bit_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \read_latency_shift_reg~1_combout ;
wire \av_readdata_pre[13]~0_combout ;


dffeas \av_readdata_pre[0] (
	.clk(clk),
	.d(av_readdata[0]),
	.asdata(q_b_0),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(read_0),
	.ena(vcc),
	.q(av_readdata_pre_0),
	.prn(vcc));
defparam \av_readdata_pre[0] .is_wysiwyg = "true";
defparam \av_readdata_pre[0] .power_up = "low";

dffeas \av_readdata_pre[16] (
	.clk(clk),
	.d(av_readdata[16]),
	.asdata(counter_reg_bit_0),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(read_0),
	.ena(vcc),
	.q(av_readdata_pre_16),
	.prn(vcc));
defparam \av_readdata_pre[16] .is_wysiwyg = "true";
defparam \av_readdata_pre[16] .power_up = "low";

dffeas \av_readdata_pre[5] (
	.clk(clk),
	.d(av_readdata[5]),
	.asdata(q_b_5),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(read_0),
	.ena(vcc),
	.q(av_readdata_pre_5),
	.prn(vcc));
defparam \av_readdata_pre[5] .is_wysiwyg = "true";
defparam \av_readdata_pre[5] .power_up = "low";

dffeas \av_readdata_pre[21] (
	.clk(clk),
	.d(av_readdata[21]),
	.asdata(counter_reg_bit_5),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(read_0),
	.ena(vcc),
	.q(av_readdata_pre_21),
	.prn(vcc));
defparam \av_readdata_pre[21] .is_wysiwyg = "true";
defparam \av_readdata_pre[21] .power_up = "low";

dffeas \av_readdata_pre[4] (
	.clk(clk),
	.d(av_readdata[5]),
	.asdata(q_b_4),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(read_0),
	.ena(vcc),
	.q(av_readdata_pre_4),
	.prn(vcc));
defparam \av_readdata_pre[4] .is_wysiwyg = "true";
defparam \av_readdata_pre[4] .power_up = "low";

dffeas \av_readdata_pre[20] (
	.clk(clk),
	.d(av_readdata[20]),
	.asdata(counter_reg_bit_4),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(read_0),
	.ena(vcc),
	.q(av_readdata_pre_20),
	.prn(vcc));
defparam \av_readdata_pre[20] .is_wysiwyg = "true";
defparam \av_readdata_pre[20] .power_up = "low";

dffeas \av_readdata_pre[6] (
	.clk(clk),
	.d(av_readdata[5]),
	.asdata(q_b_6),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(read_0),
	.ena(vcc),
	.q(av_readdata_pre_6),
	.prn(vcc));
defparam \av_readdata_pre[6] .is_wysiwyg = "true";
defparam \av_readdata_pre[6] .power_up = "low";

dffeas \av_readdata_pre[22] (
	.clk(clk),
	.d(av_readdata[22]),
	.asdata(b_full),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(read_0),
	.ena(vcc),
	.q(av_readdata_pre_22),
	.prn(vcc));
defparam \av_readdata_pre[22] .is_wysiwyg = "true";
defparam \av_readdata_pre[22] .power_up = "low";

dffeas \av_readdata_pre[7] (
	.clk(clk),
	.d(av_readdata[5]),
	.asdata(q_b_7),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(read_0),
	.ena(vcc),
	.q(av_readdata_pre_7),
	.prn(vcc));
defparam \av_readdata_pre[7] .is_wysiwyg = "true";
defparam \av_readdata_pre[7] .power_up = "low";

dffeas \av_readdata_pre[3] (
	.clk(clk),
	.d(av_readdata[5]),
	.asdata(q_b_3),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(read_0),
	.ena(vcc),
	.q(av_readdata_pre_3),
	.prn(vcc));
defparam \av_readdata_pre[3] .is_wysiwyg = "true";
defparam \av_readdata_pre[3] .power_up = "low";

dffeas \av_readdata_pre[19] (
	.clk(clk),
	.d(av_readdata[19]),
	.asdata(counter_reg_bit_3),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(read_0),
	.ena(vcc),
	.q(av_readdata_pre_19),
	.prn(vcc));
defparam \av_readdata_pre[19] .is_wysiwyg = "true";
defparam \av_readdata_pre[19] .power_up = "low";

dffeas \av_readdata_pre[2] (
	.clk(clk),
	.d(av_readdata[5]),
	.asdata(q_b_2),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(read_0),
	.ena(vcc),
	.q(av_readdata_pre_2),
	.prn(vcc));
defparam \av_readdata_pre[2] .is_wysiwyg = "true";
defparam \av_readdata_pre[2] .power_up = "low";

dffeas \av_readdata_pre[18] (
	.clk(clk),
	.d(av_readdata[18]),
	.asdata(counter_reg_bit_2),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(read_0),
	.ena(vcc),
	.q(av_readdata_pre_18),
	.prn(vcc));
defparam \av_readdata_pre[18] .is_wysiwyg = "true";
defparam \av_readdata_pre[18] .power_up = "low";

dffeas \av_readdata_pre[1] (
	.clk(clk),
	.d(av_readdata[1]),
	.asdata(q_b_1),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(read_0),
	.ena(vcc),
	.q(av_readdata_pre_1),
	.prn(vcc));
defparam \av_readdata_pre[1] .is_wysiwyg = "true";
defparam \av_readdata_pre[1] .power_up = "low";

dffeas \av_readdata_pre[17] (
	.clk(clk),
	.d(av_readdata[17]),
	.asdata(counter_reg_bit_1),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(read_0),
	.ena(vcc),
	.q(av_readdata_pre_17),
	.prn(vcc));
defparam \av_readdata_pre[17] .is_wysiwyg = "true";
defparam \av_readdata_pre[17] .power_up = "low";

dffeas \read_latency_shift_reg[0] (
	.clk(clk),
	.d(\read_latency_shift_reg~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_latency_shift_reg_0),
	.prn(vcc));
defparam \read_latency_shift_reg[0] .is_wysiwyg = "true";
defparam \read_latency_shift_reg[0] .power_up = "low";

cyclonev_lcell_comb \read_latency_shift_reg~0 (
	.dataa(!clr_break_line),
	.datab(!mem_used_1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(read_latency_shift_reg),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_latency_shift_reg~0 .extended_lut = "off";
defparam \read_latency_shift_reg~0 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \read_latency_shift_reg~0 .shared_arith = "off";

dffeas \av_readdata_pre[8] (
	.clk(clk),
	.d(av_readdata[8]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_8),
	.prn(vcc));
defparam \av_readdata_pre[8] .is_wysiwyg = "true";
defparam \av_readdata_pre[8] .power_up = "low";

dffeas \av_readdata_pre[13] (
	.clk(clk),
	.d(\av_readdata_pre[13]~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_13),
	.prn(vcc));
defparam \av_readdata_pre[13] .is_wysiwyg = "true";
defparam \av_readdata_pre[13] .power_up = "low";

dffeas \av_readdata_pre[12] (
	.clk(clk),
	.d(av_readdata[12]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_12),
	.prn(vcc));
defparam \av_readdata_pre[12] .is_wysiwyg = "true";
defparam \av_readdata_pre[12] .power_up = "low";

dffeas \av_readdata_pre[14] (
	.clk(clk),
	.d(av_readdata[14]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_14),
	.prn(vcc));
defparam \av_readdata_pre[14] .is_wysiwyg = "true";
defparam \av_readdata_pre[14] .power_up = "low";

dffeas \av_readdata_pre[15] (
	.clk(clk),
	.d(av_readdata[15]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_15),
	.prn(vcc));
defparam \av_readdata_pre[15] .is_wysiwyg = "true";
defparam \av_readdata_pre[15] .power_up = "low";

dffeas \av_readdata_pre[10] (
	.clk(clk),
	.d(av_readdata[10]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_10),
	.prn(vcc));
defparam \av_readdata_pre[10] .is_wysiwyg = "true";
defparam \av_readdata_pre[10] .power_up = "low";

dffeas \av_readdata_pre[9] (
	.clk(clk),
	.d(av_readdata[9]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_9),
	.prn(vcc));
defparam \av_readdata_pre[9] .is_wysiwyg = "true";
defparam \av_readdata_pre[9] .power_up = "low";

cyclonev_lcell_comb \read_latency_shift_reg~1 (
	.dataa(!av_waitrequest),
	.datab(!Equal6),
	.datac(!uav_read),
	.datad(!read_latency_shift_reg),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_latency_shift_reg~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_latency_shift_reg~1 .extended_lut = "off";
defparam \read_latency_shift_reg~1 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \read_latency_shift_reg~1 .shared_arith = "off";

cyclonev_lcell_comb \av_readdata_pre[13]~0 (
	.dataa(!b_full1),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_readdata_pre[13]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_readdata_pre[13]~0 .extended_lut = "off";
defparam \av_readdata_pre[13]~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \av_readdata_pre[13]~0 .shared_arith = "off";

endmodule

module processor_altera_merlin_slave_translator_2 (
	reset,
	clr_break_line,
	d_write,
	mem_used_1,
	Equal4,
	wait_latency_counter_1,
	wait_latency_counter_0,
	read_latency_shift_reg_0,
	av_waitrequest_generated,
	mem_used_11,
	src2_valid,
	av_readdata_pre_0,
	av_readdata_pre_8,
	av_readdata_pre_5,
	av_readdata_pre_4,
	av_readdata_pre_6,
	av_readdata_pre_7,
	av_readdata_pre_9,
	av_readdata_pre_3,
	av_readdata_pre_2,
	av_readdata_pre_1,
	av_readdata,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset;
input 	clr_break_line;
input 	d_write;
input 	mem_used_1;
input 	Equal4;
output 	wait_latency_counter_1;
output 	wait_latency_counter_0;
output 	read_latency_shift_reg_0;
output 	av_waitrequest_generated;
input 	mem_used_11;
input 	src2_valid;
output 	av_readdata_pre_0;
output 	av_readdata_pre_8;
output 	av_readdata_pre_5;
output 	av_readdata_pre_4;
output 	av_readdata_pre_6;
output 	av_readdata_pre_7;
output 	av_readdata_pre_9;
output 	av_readdata_pre_3;
output 	av_readdata_pre_2;
output 	av_readdata_pre_1;
input 	[31:0] av_readdata;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \wait_latency_counter[1]~0_combout ;
wire \wait_latency_counter~1_combout ;
wire \wait_latency_counter~2_combout ;
wire \read_latency_shift_reg~0_combout ;


dffeas \wait_latency_counter[1] (
	.clk(clk),
	.d(\wait_latency_counter~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wait_latency_counter_1),
	.prn(vcc));
defparam \wait_latency_counter[1] .is_wysiwyg = "true";
defparam \wait_latency_counter[1] .power_up = "low";

dffeas \wait_latency_counter[0] (
	.clk(clk),
	.d(\wait_latency_counter~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wait_latency_counter_0),
	.prn(vcc));
defparam \wait_latency_counter[0] .is_wysiwyg = "true";
defparam \wait_latency_counter[0] .power_up = "low";

dffeas \read_latency_shift_reg[0] (
	.clk(clk),
	.d(\read_latency_shift_reg~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_latency_shift_reg_0),
	.prn(vcc));
defparam \read_latency_shift_reg[0] .is_wysiwyg = "true";
defparam \read_latency_shift_reg[0] .power_up = "low";

cyclonev_lcell_comb \av_waitrequest_generated~0 (
	.dataa(!wait_latency_counter_0),
	.datab(!clr_break_line),
	.datac(!d_write),
	.datad(!mem_used_1),
	.datae(!Equal4),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(av_waitrequest_generated),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_waitrequest_generated~0 .extended_lut = "off";
defparam \av_waitrequest_generated~0 .lut_mask = 64'h9669699696696996;
defparam \av_waitrequest_generated~0 .shared_arith = "off";

dffeas \av_readdata_pre[0] (
	.clk(clk),
	.d(av_readdata[0]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_0),
	.prn(vcc));
defparam \av_readdata_pre[0] .is_wysiwyg = "true";
defparam \av_readdata_pre[0] .power_up = "low";

dffeas \av_readdata_pre[8] (
	.clk(clk),
	.d(av_readdata[8]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_8),
	.prn(vcc));
defparam \av_readdata_pre[8] .is_wysiwyg = "true";
defparam \av_readdata_pre[8] .power_up = "low";

dffeas \av_readdata_pre[5] (
	.clk(clk),
	.d(av_readdata[5]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_5),
	.prn(vcc));
defparam \av_readdata_pre[5] .is_wysiwyg = "true";
defparam \av_readdata_pre[5] .power_up = "low";

dffeas \av_readdata_pre[4] (
	.clk(clk),
	.d(av_readdata[4]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_4),
	.prn(vcc));
defparam \av_readdata_pre[4] .is_wysiwyg = "true";
defparam \av_readdata_pre[4] .power_up = "low";

dffeas \av_readdata_pre[6] (
	.clk(clk),
	.d(av_readdata[6]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_6),
	.prn(vcc));
defparam \av_readdata_pre[6] .is_wysiwyg = "true";
defparam \av_readdata_pre[6] .power_up = "low";

dffeas \av_readdata_pre[7] (
	.clk(clk),
	.d(av_readdata[7]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_7),
	.prn(vcc));
defparam \av_readdata_pre[7] .is_wysiwyg = "true";
defparam \av_readdata_pre[7] .power_up = "low";

dffeas \av_readdata_pre[9] (
	.clk(clk),
	.d(av_readdata[9]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_9),
	.prn(vcc));
defparam \av_readdata_pre[9] .is_wysiwyg = "true";
defparam \av_readdata_pre[9] .power_up = "low";

dffeas \av_readdata_pre[3] (
	.clk(clk),
	.d(av_readdata[3]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_3),
	.prn(vcc));
defparam \av_readdata_pre[3] .is_wysiwyg = "true";
defparam \av_readdata_pre[3] .power_up = "low";

dffeas \av_readdata_pre[2] (
	.clk(clk),
	.d(av_readdata[2]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_2),
	.prn(vcc));
defparam \av_readdata_pre[2] .is_wysiwyg = "true";
defparam \av_readdata_pre[2] .power_up = "low";

dffeas \av_readdata_pre[1] (
	.clk(clk),
	.d(av_readdata[1]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_1),
	.prn(vcc));
defparam \av_readdata_pre[1] .is_wysiwyg = "true";
defparam \av_readdata_pre[1] .power_up = "low";

cyclonev_lcell_comb \wait_latency_counter[1]~0 (
	.dataa(!wait_latency_counter_1),
	.datab(!mem_used_1),
	.datac(!Equal4),
	.datad(!av_waitrequest_generated),
	.datae(!src2_valid),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_latency_counter[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_latency_counter[1]~0 .extended_lut = "off";
defparam \wait_latency_counter[1]~0 .lut_mask = 64'hFFDFFFFFFFDFFFFF;
defparam \wait_latency_counter[1]~0 .shared_arith = "off";

cyclonev_lcell_comb \wait_latency_counter~1 (
	.dataa(!wait_latency_counter_1),
	.datab(!wait_latency_counter_0),
	.datac(!\wait_latency_counter[1]~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_latency_counter~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_latency_counter~1 .extended_lut = "off";
defparam \wait_latency_counter~1 .lut_mask = 64'h6F6F6F6F6F6F6F6F;
defparam \wait_latency_counter~1 .shared_arith = "off";

cyclonev_lcell_comb \wait_latency_counter~2 (
	.dataa(!wait_latency_counter_0),
	.datab(!\wait_latency_counter[1]~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_latency_counter~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_latency_counter~2 .extended_lut = "off";
defparam \wait_latency_counter~2 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \wait_latency_counter~2 .shared_arith = "off";

cyclonev_lcell_comb \read_latency_shift_reg~0 (
	.dataa(!mem_used_1),
	.datab(!mem_used_11),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_latency_shift_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_latency_shift_reg~0 .extended_lut = "off";
defparam \read_latency_shift_reg~0 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \read_latency_shift_reg~0 .shared_arith = "off";

endmodule

module processor_altera_merlin_slave_translator_3 (
	reset,
	clr_break_line,
	read_latency_shift_reg_0,
	mem_used_1,
	read_latency_shift_reg,
	rf_source_valid,
	read_latency_shift_reg1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset;
input 	clr_break_line;
output 	read_latency_shift_reg_0;
input 	mem_used_1;
output 	read_latency_shift_reg;
input 	rf_source_valid;
output 	read_latency_shift_reg1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \read_latency_shift_reg[0] (
	.clk(clk),
	.d(read_latency_shift_reg1),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_latency_shift_reg_0),
	.prn(vcc));
defparam \read_latency_shift_reg[0] .is_wysiwyg = "true";
defparam \read_latency_shift_reg[0] .power_up = "low";

cyclonev_lcell_comb \read_latency_shift_reg~0 (
	.dataa(!clr_break_line),
	.datab(!mem_used_1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(read_latency_shift_reg),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_latency_shift_reg~0 .extended_lut = "off";
defparam \read_latency_shift_reg~0 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \read_latency_shift_reg~0 .shared_arith = "off";

cyclonev_lcell_comb \read_latency_shift_reg~1 (
	.dataa(!read_latency_shift_reg),
	.datab(!rf_source_valid),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(read_latency_shift_reg1),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_latency_shift_reg~1 .extended_lut = "off";
defparam \read_latency_shift_reg~1 .lut_mask = 64'h7777777777777777;
defparam \read_latency_shift_reg~1 .shared_arith = "off";

endmodule

module processor_altera_merlin_slave_translator_4 (
	reset,
	d_write,
	read_latency_shift_reg_0,
	sink_ready,
	wait_latency_counter_1,
	wait_latency_counter_0,
	sink_ready1,
	uav_read,
	av_readdata_pre_0,
	av_readdata_pre_8,
	av_readdata_pre_5,
	av_readdata_pre_4,
	av_readdata_pre_6,
	av_readdata_pre_7,
	av_readdata_pre_9,
	av_readdata_pre_3,
	av_readdata_pre_2,
	av_readdata_pre_1,
	av_readdata,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset;
input 	d_write;
output 	read_latency_shift_reg_0;
input 	sink_ready;
output 	wait_latency_counter_1;
output 	wait_latency_counter_0;
input 	sink_ready1;
input 	uav_read;
output 	av_readdata_pre_0;
output 	av_readdata_pre_8;
output 	av_readdata_pre_5;
output 	av_readdata_pre_4;
output 	av_readdata_pre_6;
output 	av_readdata_pre_7;
output 	av_readdata_pre_9;
output 	av_readdata_pre_3;
output 	av_readdata_pre_2;
output 	av_readdata_pre_1;
input 	[31:0] av_readdata;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \wait_latency_counter~0_combout ;
wire \wait_latency_counter~1_combout ;


dffeas \read_latency_shift_reg[0] (
	.clk(clk),
	.d(sink_ready1),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_latency_shift_reg_0),
	.prn(vcc));
defparam \read_latency_shift_reg[0] .is_wysiwyg = "true";
defparam \read_latency_shift_reg[0] .power_up = "low";

dffeas \wait_latency_counter[1] (
	.clk(clk),
	.d(\wait_latency_counter~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wait_latency_counter_1),
	.prn(vcc));
defparam \wait_latency_counter[1] .is_wysiwyg = "true";
defparam \wait_latency_counter[1] .power_up = "low";

dffeas \wait_latency_counter[0] (
	.clk(clk),
	.d(\wait_latency_counter~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wait_latency_counter_0),
	.prn(vcc));
defparam \wait_latency_counter[0] .is_wysiwyg = "true";
defparam \wait_latency_counter[0] .power_up = "low";

dffeas \av_readdata_pre[0] (
	.clk(clk),
	.d(av_readdata[0]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_0),
	.prn(vcc));
defparam \av_readdata_pre[0] .is_wysiwyg = "true";
defparam \av_readdata_pre[0] .power_up = "low";

dffeas \av_readdata_pre[8] (
	.clk(clk),
	.d(av_readdata[8]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_8),
	.prn(vcc));
defparam \av_readdata_pre[8] .is_wysiwyg = "true";
defparam \av_readdata_pre[8] .power_up = "low";

dffeas \av_readdata_pre[5] (
	.clk(clk),
	.d(av_readdata[5]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_5),
	.prn(vcc));
defparam \av_readdata_pre[5] .is_wysiwyg = "true";
defparam \av_readdata_pre[5] .power_up = "low";

dffeas \av_readdata_pre[4] (
	.clk(clk),
	.d(av_readdata[4]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_4),
	.prn(vcc));
defparam \av_readdata_pre[4] .is_wysiwyg = "true";
defparam \av_readdata_pre[4] .power_up = "low";

dffeas \av_readdata_pre[6] (
	.clk(clk),
	.d(av_readdata[6]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_6),
	.prn(vcc));
defparam \av_readdata_pre[6] .is_wysiwyg = "true";
defparam \av_readdata_pre[6] .power_up = "low";

dffeas \av_readdata_pre[7] (
	.clk(clk),
	.d(av_readdata[7]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_7),
	.prn(vcc));
defparam \av_readdata_pre[7] .is_wysiwyg = "true";
defparam \av_readdata_pre[7] .power_up = "low";

dffeas \av_readdata_pre[9] (
	.clk(clk),
	.d(av_readdata[9]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_9),
	.prn(vcc));
defparam \av_readdata_pre[9] .is_wysiwyg = "true";
defparam \av_readdata_pre[9] .power_up = "low";

dffeas \av_readdata_pre[3] (
	.clk(clk),
	.d(av_readdata[3]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_3),
	.prn(vcc));
defparam \av_readdata_pre[3] .is_wysiwyg = "true";
defparam \av_readdata_pre[3] .power_up = "low";

dffeas \av_readdata_pre[2] (
	.clk(clk),
	.d(av_readdata[2]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_2),
	.prn(vcc));
defparam \av_readdata_pre[2] .is_wysiwyg = "true";
defparam \av_readdata_pre[2] .power_up = "low";

dffeas \av_readdata_pre[1] (
	.clk(clk),
	.d(av_readdata[1]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_1),
	.prn(vcc));
defparam \av_readdata_pre[1] .is_wysiwyg = "true";
defparam \av_readdata_pre[1] .power_up = "low";

cyclonev_lcell_comb \wait_latency_counter~0 (
	.dataa(!d_write),
	.datab(!uav_read),
	.datac(!sink_ready),
	.datad(!wait_latency_counter_1),
	.datae(!wait_latency_counter_0),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_latency_counter~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_latency_counter~0 .extended_lut = "off";
defparam \wait_latency_counter~0 .lut_mask = 64'h7FFFFF7F7FFFFF7F;
defparam \wait_latency_counter~0 .shared_arith = "off";

cyclonev_lcell_comb \wait_latency_counter~1 (
	.dataa(!d_write),
	.datab(!uav_read),
	.datac(!sink_ready),
	.datad(!wait_latency_counter_1),
	.datae(!wait_latency_counter_0),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_latency_counter~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_latency_counter~1 .extended_lut = "off";
defparam \wait_latency_counter~1 .lut_mask = 64'hBFFF1FFFBFFF1FFF;
defparam \wait_latency_counter~1 .shared_arith = "off";

endmodule

module processor_altera_merlin_slave_translator_5 (
	reset,
	d_write,
	read_latency_shift_reg_0,
	wait_latency_counter_1,
	wait_latency_counter_0,
	uav_read,
	period_l_wr_strobe,
	mem_used_1,
	read_latency_shift_reg,
	av_readdata_pre_0,
	av_readdata_pre_8,
	av_readdata_pre_5,
	av_readdata_pre_13,
	av_readdata_pre_4,
	av_readdata_pre_12,
	av_readdata_pre_6,
	av_readdata_pre_14,
	av_readdata_pre_7,
	av_readdata_pre_15,
	av_readdata_pre_11,
	av_readdata_pre_10,
	av_readdata_pre_9,
	av_readdata_pre_3,
	av_readdata_pre_2,
	av_readdata_pre_1,
	av_readdata,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset;
input 	d_write;
output 	read_latency_shift_reg_0;
output 	wait_latency_counter_1;
output 	wait_latency_counter_0;
input 	uav_read;
input 	period_l_wr_strobe;
input 	mem_used_1;
output 	read_latency_shift_reg;
output 	av_readdata_pre_0;
output 	av_readdata_pre_8;
output 	av_readdata_pre_5;
output 	av_readdata_pre_13;
output 	av_readdata_pre_4;
output 	av_readdata_pre_12;
output 	av_readdata_pre_6;
output 	av_readdata_pre_14;
output 	av_readdata_pre_7;
output 	av_readdata_pre_15;
output 	av_readdata_pre_11;
output 	av_readdata_pre_10;
output 	av_readdata_pre_9;
output 	av_readdata_pre_3;
output 	av_readdata_pre_2;
output 	av_readdata_pre_1;
input 	[31:0] av_readdata;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \wait_latency_counter~0_combout ;
wire \wait_latency_counter~1_combout ;


dffeas \read_latency_shift_reg[0] (
	.clk(clk),
	.d(read_latency_shift_reg),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_latency_shift_reg_0),
	.prn(vcc));
defparam \read_latency_shift_reg[0] .is_wysiwyg = "true";
defparam \read_latency_shift_reg[0] .power_up = "low";

dffeas \wait_latency_counter[1] (
	.clk(clk),
	.d(\wait_latency_counter~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wait_latency_counter_1),
	.prn(vcc));
defparam \wait_latency_counter[1] .is_wysiwyg = "true";
defparam \wait_latency_counter[1] .power_up = "low";

dffeas \wait_latency_counter[0] (
	.clk(clk),
	.d(\wait_latency_counter~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wait_latency_counter_0),
	.prn(vcc));
defparam \wait_latency_counter[0] .is_wysiwyg = "true";
defparam \wait_latency_counter[0] .power_up = "low";

cyclonev_lcell_comb \read_latency_shift_reg~0 (
	.dataa(!period_l_wr_strobe),
	.datab(!mem_used_1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(read_latency_shift_reg),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_latency_shift_reg~0 .extended_lut = "off";
defparam \read_latency_shift_reg~0 .lut_mask = 64'h7777777777777777;
defparam \read_latency_shift_reg~0 .shared_arith = "off";

dffeas \av_readdata_pre[0] (
	.clk(clk),
	.d(av_readdata[0]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_0),
	.prn(vcc));
defparam \av_readdata_pre[0] .is_wysiwyg = "true";
defparam \av_readdata_pre[0] .power_up = "low";

dffeas \av_readdata_pre[8] (
	.clk(clk),
	.d(av_readdata[8]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_8),
	.prn(vcc));
defparam \av_readdata_pre[8] .is_wysiwyg = "true";
defparam \av_readdata_pre[8] .power_up = "low";

dffeas \av_readdata_pre[5] (
	.clk(clk),
	.d(av_readdata[5]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_5),
	.prn(vcc));
defparam \av_readdata_pre[5] .is_wysiwyg = "true";
defparam \av_readdata_pre[5] .power_up = "low";

dffeas \av_readdata_pre[13] (
	.clk(clk),
	.d(av_readdata[13]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_13),
	.prn(vcc));
defparam \av_readdata_pre[13] .is_wysiwyg = "true";
defparam \av_readdata_pre[13] .power_up = "low";

dffeas \av_readdata_pre[4] (
	.clk(clk),
	.d(av_readdata[4]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_4),
	.prn(vcc));
defparam \av_readdata_pre[4] .is_wysiwyg = "true";
defparam \av_readdata_pre[4] .power_up = "low";

dffeas \av_readdata_pre[12] (
	.clk(clk),
	.d(av_readdata[12]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_12),
	.prn(vcc));
defparam \av_readdata_pre[12] .is_wysiwyg = "true";
defparam \av_readdata_pre[12] .power_up = "low";

dffeas \av_readdata_pre[6] (
	.clk(clk),
	.d(av_readdata[6]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_6),
	.prn(vcc));
defparam \av_readdata_pre[6] .is_wysiwyg = "true";
defparam \av_readdata_pre[6] .power_up = "low";

dffeas \av_readdata_pre[14] (
	.clk(clk),
	.d(av_readdata[14]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_14),
	.prn(vcc));
defparam \av_readdata_pre[14] .is_wysiwyg = "true";
defparam \av_readdata_pre[14] .power_up = "low";

dffeas \av_readdata_pre[7] (
	.clk(clk),
	.d(av_readdata[7]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_7),
	.prn(vcc));
defparam \av_readdata_pre[7] .is_wysiwyg = "true";
defparam \av_readdata_pre[7] .power_up = "low";

dffeas \av_readdata_pre[15] (
	.clk(clk),
	.d(av_readdata[15]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_15),
	.prn(vcc));
defparam \av_readdata_pre[15] .is_wysiwyg = "true";
defparam \av_readdata_pre[15] .power_up = "low";

dffeas \av_readdata_pre[11] (
	.clk(clk),
	.d(av_readdata[11]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_11),
	.prn(vcc));
defparam \av_readdata_pre[11] .is_wysiwyg = "true";
defparam \av_readdata_pre[11] .power_up = "low";

dffeas \av_readdata_pre[10] (
	.clk(clk),
	.d(av_readdata[10]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_10),
	.prn(vcc));
defparam \av_readdata_pre[10] .is_wysiwyg = "true";
defparam \av_readdata_pre[10] .power_up = "low";

dffeas \av_readdata_pre[9] (
	.clk(clk),
	.d(av_readdata[9]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_9),
	.prn(vcc));
defparam \av_readdata_pre[9] .is_wysiwyg = "true";
defparam \av_readdata_pre[9] .power_up = "low";

dffeas \av_readdata_pre[3] (
	.clk(clk),
	.d(av_readdata[3]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_3),
	.prn(vcc));
defparam \av_readdata_pre[3] .is_wysiwyg = "true";
defparam \av_readdata_pre[3] .power_up = "low";

dffeas \av_readdata_pre[2] (
	.clk(clk),
	.d(av_readdata[2]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_2),
	.prn(vcc));
defparam \av_readdata_pre[2] .is_wysiwyg = "true";
defparam \av_readdata_pre[2] .power_up = "low";

dffeas \av_readdata_pre[1] (
	.clk(clk),
	.d(av_readdata[1]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_1),
	.prn(vcc));
defparam \av_readdata_pre[1] .is_wysiwyg = "true";
defparam \av_readdata_pre[1] .power_up = "low";

cyclonev_lcell_comb \wait_latency_counter~0 (
	.dataa(!d_write),
	.datab(!uav_read),
	.datac(!wait_latency_counter_1),
	.datad(!wait_latency_counter_0),
	.datae(!period_l_wr_strobe),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_latency_counter~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_latency_counter~0 .extended_lut = "off";
defparam \wait_latency_counter~0 .lut_mask = 64'h7FF7FFFF7FF7FFFF;
defparam \wait_latency_counter~0 .shared_arith = "off";

cyclonev_lcell_comb \wait_latency_counter~1 (
	.dataa(!d_write),
	.datab(!uav_read),
	.datac(!wait_latency_counter_1),
	.datad(!wait_latency_counter_0),
	.datae(!period_l_wr_strobe),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_latency_counter~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_latency_counter~1 .extended_lut = "off";
defparam \wait_latency_counter~1 .lut_mask = 64'hBF1FFFFFBF1FFFFF;
defparam \wait_latency_counter~1 .shared_arith = "off";

endmodule

module processor_altera_merlin_slave_translator_6 (
	reset,
	d_write,
	av_readdata,
	read_latency_shift_reg_0,
	sink_ready,
	wait_latency_counter_1,
	wait_latency_counter_0,
	sink_ready1,
	uav_read,
	av_readdata_pre_30,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset;
input 	d_write;
input 	[31:0] av_readdata;
output 	read_latency_shift_reg_0;
input 	sink_ready;
output 	wait_latency_counter_1;
output 	wait_latency_counter_0;
input 	sink_ready1;
input 	uav_read;
output 	av_readdata_pre_30;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \wait_latency_counter~0_combout ;
wire \wait_latency_counter~1_combout ;


dffeas \read_latency_shift_reg[0] (
	.clk(clk),
	.d(sink_ready1),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_latency_shift_reg_0),
	.prn(vcc));
defparam \read_latency_shift_reg[0] .is_wysiwyg = "true";
defparam \read_latency_shift_reg[0] .power_up = "low";

dffeas \wait_latency_counter[1] (
	.clk(clk),
	.d(\wait_latency_counter~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wait_latency_counter_1),
	.prn(vcc));
defparam \wait_latency_counter[1] .is_wysiwyg = "true";
defparam \wait_latency_counter[1] .power_up = "low";

dffeas \wait_latency_counter[0] (
	.clk(clk),
	.d(\wait_latency_counter~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wait_latency_counter_0),
	.prn(vcc));
defparam \wait_latency_counter[0] .is_wysiwyg = "true";
defparam \wait_latency_counter[0] .power_up = "low";

dffeas \av_readdata_pre[30] (
	.clk(clk),
	.d(av_readdata[30]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_30),
	.prn(vcc));
defparam \av_readdata_pre[30] .is_wysiwyg = "true";
defparam \av_readdata_pre[30] .power_up = "low";

cyclonev_lcell_comb \wait_latency_counter~0 (
	.dataa(!d_write),
	.datab(!uav_read),
	.datac(!sink_ready),
	.datad(!wait_latency_counter_1),
	.datae(!wait_latency_counter_0),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_latency_counter~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_latency_counter~0 .extended_lut = "off";
defparam \wait_latency_counter~0 .lut_mask = 64'h7FFFFF7F7FFFFF7F;
defparam \wait_latency_counter~0 .shared_arith = "off";

cyclonev_lcell_comb \wait_latency_counter~1 (
	.dataa(!d_write),
	.datab(!uav_read),
	.datac(!sink_ready),
	.datad(!wait_latency_counter_1),
	.datae(!wait_latency_counter_0),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_latency_counter~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_latency_counter~1 .extended_lut = "off";
defparam \wait_latency_counter~1 .lut_mask = 64'hBFFF1FFFBFFF1FFF;
defparam \wait_latency_counter~1 .shared_arith = "off";

endmodule

module processor_altera_merlin_traffic_limiter (
	reset,
	clr_break_line,
	i_read,
	last_channel_0,
	has_pending_responses1,
	cmd_sink_channel,
	last_dest_id_1,
	WideOr0,
	nonposted_cmd_accepted1,
	src1_valid,
	src1_valid1,
	mem_61_0,
	mem_61_01,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset;
input 	clr_break_line;
input 	i_read;
output 	last_channel_0;
output 	has_pending_responses1;
input 	[6:0] cmd_sink_channel;
output 	last_dest_id_1;
input 	WideOr0;
output 	nonposted_cmd_accepted1;
input 	src1_valid;
input 	src1_valid1;
input 	mem_61_0;
input 	mem_61_01;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \save_dest_id~0_combout ;
wire \response_sink_accepted~0_combout ;
wire \pending_response_count[0]~0_combout ;
wire \pending_response_count[0]~q ;
wire \has_pending_responses~0_combout ;
wire \last_dest_id[1]~0_combout ;


dffeas \last_channel[0] (
	.clk(clk),
	.d(cmd_sink_channel[0]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\save_dest_id~0_combout ),
	.q(last_channel_0),
	.prn(vcc));
defparam \last_channel[0] .is_wysiwyg = "true";
defparam \last_channel[0] .power_up = "low";

dffeas has_pending_responses(
	.clk(clk),
	.d(\has_pending_responses~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(has_pending_responses1),
	.prn(vcc));
defparam has_pending_responses.is_wysiwyg = "true";
defparam has_pending_responses.power_up = "low";

dffeas \last_dest_id[1] (
	.clk(clk),
	.d(\last_dest_id[1]~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\save_dest_id~0_combout ),
	.q(last_dest_id_1),
	.prn(vcc));
defparam \last_dest_id[1] .is_wysiwyg = "true";
defparam \last_dest_id[1] .power_up = "low";

cyclonev_lcell_comb nonposted_cmd_accepted(
	.dataa(!\save_dest_id~0_combout ),
	.datab(!WideOr0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(nonposted_cmd_accepted1),
	.sumout(),
	.cout(),
	.shareout());
defparam nonposted_cmd_accepted.extended_lut = "off";
defparam nonposted_cmd_accepted.lut_mask = 64'h7777777777777777;
defparam nonposted_cmd_accepted.shared_arith = "off";

cyclonev_lcell_comb \save_dest_id~0 (
	.dataa(!clr_break_line),
	.datab(!has_pending_responses1),
	.datac(!i_read),
	.datad(!cmd_sink_channel[0]),
	.datae(!last_dest_id_1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\save_dest_id~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \save_dest_id~0 .extended_lut = "off";
defparam \save_dest_id~0 .lut_mask = 64'hDFFFFFDFDFFFFFDF;
defparam \save_dest_id~0 .shared_arith = "off";

cyclonev_lcell_comb \response_sink_accepted~0 (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!mem_61_0),
	.datad(!mem_61_01),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\response_sink_accepted~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \response_sink_accepted~0 .extended_lut = "off";
defparam \response_sink_accepted~0 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \response_sink_accepted~0 .shared_arith = "off";

cyclonev_lcell_comb \pending_response_count[0]~0 (
	.dataa(!nonposted_cmd_accepted1),
	.datab(!\pending_response_count[0]~q ),
	.datac(!\response_sink_accepted~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pending_response_count[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pending_response_count[0]~0 .extended_lut = "off";
defparam \pending_response_count[0]~0 .lut_mask = 64'h9696969696969696;
defparam \pending_response_count[0]~0 .shared_arith = "off";

dffeas \pending_response_count[0] (
	.clk(clk),
	.d(\pending_response_count[0]~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\pending_response_count[0]~q ),
	.prn(vcc));
defparam \pending_response_count[0] .is_wysiwyg = "true";
defparam \pending_response_count[0] .power_up = "low";

cyclonev_lcell_comb \has_pending_responses~0 (
	.dataa(!has_pending_responses1),
	.datab(!nonposted_cmd_accepted1),
	.datac(!\pending_response_count[0]~q ),
	.datad(!\response_sink_accepted~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\has_pending_responses~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \has_pending_responses~0 .extended_lut = "off";
defparam \has_pending_responses~0 .lut_mask = 64'hFFF7FFF7FFF7FFF7;
defparam \has_pending_responses~0 .shared_arith = "off";

cyclonev_lcell_comb \last_dest_id[1]~0 (
	.dataa(!cmd_sink_channel[0]),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\last_dest_id[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_dest_id[1]~0 .extended_lut = "off";
defparam \last_dest_id[1]~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \last_dest_id[1]~0 .shared_arith = "off";

endmodule

module processor_processor_mm_interconnect_0_cmd_demux (
	clr_break_line,
	d_write,
	Equal1,
	Equal2,
	Equal4,
	d_read,
	mem_used_1,
	read_accepted,
	always1,
	always11,
	sink_ready,
	wait_latency_counter_1,
	wait_latency_counter_0,
	sink_ready1,
	mem_used_11,
	always12,
	sink_ready2,
	wait_latency_counter_11,
	wait_latency_counter_01,
	sink_ready3,
	Equal21,
	mem_used_12,
	av_waitrequest,
	Equal6,
	sink_ready4,
	saved_grant_0,
	write,
	saved_grant_01,
	read_latency_shift_reg,
	Equal11,
	WideOr0,
	src2_valid,
	src2_valid1,
	src2_valid2,
	src3_valid,
	sink_ready5,
	sink_ready6,
	sink_ready7,
	sink_ready8)/* synthesis synthesis_greybox=1 */;
input 	clr_break_line;
input 	d_write;
input 	Equal1;
input 	Equal2;
input 	Equal4;
input 	d_read;
input 	mem_used_1;
input 	read_accepted;
input 	always1;
input 	always11;
output 	sink_ready;
input 	wait_latency_counter_1;
input 	wait_latency_counter_0;
output 	sink_ready1;
input 	mem_used_11;
input 	always12;
output 	sink_ready2;
input 	wait_latency_counter_11;
input 	wait_latency_counter_01;
output 	sink_ready3;
input 	Equal21;
input 	mem_used_12;
input 	av_waitrequest;
input 	Equal6;
output 	sink_ready4;
input 	saved_grant_0;
input 	write;
input 	saved_grant_01;
input 	read_latency_shift_reg;
input 	Equal11;
output 	WideOr0;
output 	src2_valid;
output 	src2_valid1;
output 	src2_valid2;
output 	src3_valid;
output 	sink_ready5;
output 	sink_ready6;
output 	sink_ready7;
output 	sink_ready8;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \sink_ready~9_combout ;
wire \sink_ready~10_combout ;


cyclonev_lcell_comb \sink_ready~0 (
	.dataa(!clr_break_line),
	.datab(!Equal1),
	.datac(!Equal2),
	.datad(!mem_used_1),
	.datae(!always1),
	.dataf(!always11),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(sink_ready),
	.sumout(),
	.cout(),
	.shareout());
defparam \sink_ready~0 .extended_lut = "off";
defparam \sink_ready~0 .lut_mask = 64'hFF7FFFFFFFFFFFFF;
defparam \sink_ready~0 .shared_arith = "off";

cyclonev_lcell_comb \sink_ready~1 (
	.dataa(!wait_latency_counter_1),
	.datab(!Equal1),
	.datac(!Equal2),
	.datad(!always1),
	.datae(!always11),
	.dataf(!\sink_ready~9_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(sink_ready1),
	.sumout(),
	.cout(),
	.shareout());
defparam \sink_ready~1 .extended_lut = "off";
defparam \sink_ready~1 .lut_mask = 64'hBFFFFFFFFFFFFFFF;
defparam \sink_ready~1 .shared_arith = "off";

cyclonev_lcell_comb \sink_ready~2 (
	.dataa(!clr_break_line),
	.datab(!Equal1),
	.datac(!Equal2),
	.datad(!always1),
	.datae(!mem_used_11),
	.dataf(!always12),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(sink_ready2),
	.sumout(),
	.cout(),
	.shareout());
defparam \sink_ready~2 .extended_lut = "off";
defparam \sink_ready~2 .lut_mask = 64'hFFFF7FFFFFFFFFFF;
defparam \sink_ready~2 .shared_arith = "off";

cyclonev_lcell_comb \sink_ready~3 (
	.dataa(!wait_latency_counter_11),
	.datab(!Equal1),
	.datac(!Equal2),
	.datad(!always1),
	.datae(!always12),
	.dataf(!\sink_ready~10_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(sink_ready3),
	.sumout(),
	.cout(),
	.shareout());
defparam \sink_ready~3 .extended_lut = "off";
defparam \sink_ready~3 .lut_mask = 64'hBFFFFFFFFFFFFFFF;
defparam \sink_ready~3 .shared_arith = "off";

cyclonev_lcell_comb \sink_ready~4 (
	.dataa(!Equal1),
	.datab(!Equal2),
	.datac(!mem_used_12),
	.datad(!av_waitrequest),
	.datae(!Equal6),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(sink_ready4),
	.sumout(),
	.cout(),
	.shareout());
defparam \sink_ready~4 .extended_lut = "off";
defparam \sink_ready~4 .lut_mask = 64'hF7FFFFFFF7FFFFFF;
defparam \sink_ready~4 .shared_arith = "off";

cyclonev_lcell_comb \WideOr0~0 (
	.dataa(!saved_grant_0),
	.datab(!write),
	.datac(!saved_grant_01),
	.datad(!read_latency_shift_reg),
	.datae(!Equal11),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(WideOr0),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr0~0 .extended_lut = "off";
defparam \WideOr0~0 .lut_mask = 64'h5FFF3FFF5FFF3FFF;
defparam \WideOr0~0 .shared_arith = "off";

cyclonev_lcell_comb \src2_valid~0 (
	.dataa(!Equal1),
	.datab(!Equal2),
	.datac(!Equal6),
	.datad(!always1),
	.datae(!always11),
	.dataf(!always12),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src2_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src2_valid~0 .extended_lut = "off";
defparam \src2_valid~0 .lut_mask = 64'h7FFFFFFFFFFFFFFF;
defparam \src2_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \src2_valid~1 (
	.dataa(!clr_break_line),
	.datab(!d_write),
	.datac(!d_read),
	.datad(!read_accepted),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src2_valid1),
	.sumout(),
	.cout(),
	.shareout());
defparam \src2_valid~1 .extended_lut = "off";
defparam \src2_valid~1 .lut_mask = 64'hFF7FFF7FFF7FFF7F;
defparam \src2_valid~1 .shared_arith = "off";

cyclonev_lcell_comb \src2_valid~2 (
	.dataa(!Equal4),
	.datab(!Equal11),
	.datac(!Equal21),
	.datad(!src2_valid),
	.datae(!src2_valid1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src2_valid2),
	.sumout(),
	.cout(),
	.shareout());
defparam \src2_valid~2 .extended_lut = "off";
defparam \src2_valid~2 .lut_mask = 64'hFFFBFFFFFFFBFFFF;
defparam \src2_valid~2 .shared_arith = "off";

cyclonev_lcell_comb \src3_valid~0 (
	.dataa(!Equal4),
	.datab(!Equal11),
	.datac(!Equal21),
	.datad(!src2_valid),
	.datae(!src2_valid1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src3_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src3_valid~0 .extended_lut = "off";
defparam \src3_valid~0 .lut_mask = 64'hFFFEFFFFFFFEFFFF;
defparam \src3_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \sink_ready~5 (
	.dataa(!clr_break_line),
	.datab(!Equal1),
	.datac(!Equal2),
	.datad(!always1),
	.datae(!always11),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(sink_ready5),
	.sumout(),
	.cout(),
	.shareout());
defparam \sink_ready~5 .extended_lut = "off";
defparam \sink_ready~5 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \sink_ready~5 .shared_arith = "off";

cyclonev_lcell_comb \sink_ready~6 (
	.dataa(!d_write),
	.datab(!sink_ready),
	.datac(!wait_latency_counter_1),
	.datad(!wait_latency_counter_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(sink_ready6),
	.sumout(),
	.cout(),
	.shareout());
defparam \sink_ready~6 .extended_lut = "off";
defparam \sink_ready~6 .lut_mask = 64'hF9F6F9F6F9F6F9F6;
defparam \sink_ready~6 .shared_arith = "off";

cyclonev_lcell_comb \sink_ready~7 (
	.dataa(!clr_break_line),
	.datab(!Equal1),
	.datac(!Equal2),
	.datad(!always1),
	.datae(!always12),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(sink_ready7),
	.sumout(),
	.cout(),
	.shareout());
defparam \sink_ready~7 .extended_lut = "off";
defparam \sink_ready~7 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \sink_ready~7 .shared_arith = "off";

cyclonev_lcell_comb \sink_ready~8 (
	.dataa(!d_write),
	.datab(!sink_ready2),
	.datac(!wait_latency_counter_11),
	.datad(!wait_latency_counter_01),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(sink_ready8),
	.sumout(),
	.cout(),
	.shareout());
defparam \sink_ready~8 .extended_lut = "off";
defparam \sink_ready~8 .lut_mask = 64'hF9F6F9F6F9F6F9F6;
defparam \sink_ready~8 .shared_arith = "off";

cyclonev_lcell_comb \sink_ready~9 (
	.dataa(!d_write),
	.datab(!wait_latency_counter_0),
	.datac(!clr_break_line),
	.datad(!mem_used_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sink_ready~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sink_ready~9 .extended_lut = "off";
defparam \sink_ready~9 .lut_mask = 64'hFF6FFF6FFF6FFF6F;
defparam \sink_ready~9 .shared_arith = "off";

cyclonev_lcell_comb \sink_ready~10 (
	.dataa(!d_write),
	.datab(!wait_latency_counter_01),
	.datac(!clr_break_line),
	.datad(!mem_used_11),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sink_ready~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sink_ready~10 .extended_lut = "off";
defparam \sink_ready~10 .lut_mask = 64'hFF6FFF6FFF6FFF6F;
defparam \sink_ready~10 .shared_arith = "off";

endmodule

module processor_processor_mm_interconnect_0_cmd_demux_001 (
	clr_break_line,
	write,
	read_latency_shift_reg,
	saved_grant_1,
	i_read,
	last_channel_0,
	has_pending_responses,
	Equal1,
	src0_valid,
	saved_grant_11,
	last_dest_id_1,
	src1_valid,
	WideOr0)/* synthesis synthesis_greybox=1 */;
input 	clr_break_line;
input 	write;
input 	read_latency_shift_reg;
input 	saved_grant_1;
input 	i_read;
input 	last_channel_0;
input 	has_pending_responses;
input 	Equal1;
output 	src0_valid;
input 	saved_grant_11;
input 	last_dest_id_1;
output 	src1_valid;
output 	WideOr0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb \src0_valid~0 (
	.dataa(!clr_break_line),
	.datab(!last_channel_0),
	.datac(!has_pending_responses),
	.datad(!i_read),
	.datae(!Equal1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src0_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src0_valid~0 .extended_lut = "off";
defparam \src0_valid~0 .lut_mask = 64'hF7FFFFFFF7FFFFFF;
defparam \src0_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \src1_valid~0 (
	.dataa(!clr_break_line),
	.datab(!has_pending_responses),
	.datac(!i_read),
	.datad(!Equal1),
	.datae(!last_dest_id_1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src1_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src1_valid~0 .extended_lut = "off";
defparam \src1_valid~0 .lut_mask = 64'hFFDFFFFFFFDFFFFF;
defparam \src1_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \WideOr0~0 (
	.dataa(!write),
	.datab(!read_latency_shift_reg),
	.datac(!saved_grant_1),
	.datad(!Equal1),
	.datae(!saved_grant_11),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(WideOr0),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr0~0 .extended_lut = "off";
defparam \WideOr0~0 .lut_mask = 64'h5F3FFFFF5F3FFFFF;
defparam \WideOr0~0 .shared_arith = "off";

endmodule

module processor_processor_mm_interconnect_0_cmd_mux_002 (
	M_st_data_8,
	M_st_data_9,
	M_st_data_16,
	M_st_data_21,
	M_st_data_13,
	M_st_data_20,
	M_st_data_12,
	M_st_data_22,
	M_st_data_14,
	M_st_data_23,
	M_st_data_15,
	M_st_data_11,
	M_st_data_10,
	M_st_data_19,
	M_st_data_18,
	M_st_data_17,
	M_st_data_0,
	r_sync_rst,
	M_alu_result_5,
	M_alu_result_4,
	M_alu_result_6,
	M_alu_result_10,
	M_alu_result_9,
	M_alu_result_8,
	M_alu_result_7,
	M_alu_result_3,
	M_alu_result_2,
	M_st_data_1,
	M_st_data_2,
	M_st_data_3,
	M_st_data_4,
	M_st_data_5,
	M_st_data_6,
	M_st_data_7,
	saved_grant_0,
	write,
	hbreak_enabled,
	src2_valid,
	saved_grant_1,
	src0_valid,
	ic_fill_line_5,
	src_data_46,
	ic_fill_line_0,
	ic_fill_line_1,
	ic_fill_line_2,
	ic_fill_line_3,
	ic_fill_line_4,
	ic_fill_ap_offset_0,
	ic_fill_ap_offset_1,
	ic_fill_ap_offset_2,
	M_mem_byte_en_0,
	M_mem_byte_en_2,
	M_mem_byte_en_1,
	M_st_data_24,
	M_mem_byte_en_3,
	src_payload,
	src_data_38,
	src_data_41,
	src_data_40,
	src_data_39,
	src_data_45,
	src_data_44,
	src_data_43,
	src_data_42,
	src_payload1,
	M_st_data_29,
	M_st_data_28,
	M_st_data_30,
	M_st_data_31,
	M_st_data_27,
	M_st_data_26,
	M_st_data_25,
	src_payload2,
	src_data_32,
	src_payload3,
	src_payload4,
	src_payload5,
	src_data_34,
	src_payload6,
	src_data_33,
	src_payload7,
	src_data_35,
	src_payload8,
	src_payload9,
	src_payload10,
	src_payload11,
	src_payload12,
	src_payload13,
	src_payload14,
	src_payload15,
	src_payload16,
	src_payload17,
	src_payload18,
	src_payload19,
	src_payload20,
	src_payload21,
	src_payload22,
	src_payload23,
	src_payload24,
	src_payload25,
	src_payload26,
	src_payload27,
	src_payload28,
	src_payload29,
	src_payload30,
	src_payload31,
	src_payload32,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	M_st_data_8;
input 	M_st_data_9;
input 	M_st_data_16;
input 	M_st_data_21;
input 	M_st_data_13;
input 	M_st_data_20;
input 	M_st_data_12;
input 	M_st_data_22;
input 	M_st_data_14;
input 	M_st_data_23;
input 	M_st_data_15;
input 	M_st_data_11;
input 	M_st_data_10;
input 	M_st_data_19;
input 	M_st_data_18;
input 	M_st_data_17;
input 	M_st_data_0;
input 	r_sync_rst;
input 	M_alu_result_5;
input 	M_alu_result_4;
input 	M_alu_result_6;
input 	M_alu_result_10;
input 	M_alu_result_9;
input 	M_alu_result_8;
input 	M_alu_result_7;
input 	M_alu_result_3;
input 	M_alu_result_2;
input 	M_st_data_1;
input 	M_st_data_2;
input 	M_st_data_3;
input 	M_st_data_4;
input 	M_st_data_5;
input 	M_st_data_6;
input 	M_st_data_7;
output 	saved_grant_0;
input 	write;
input 	hbreak_enabled;
input 	src2_valid;
output 	saved_grant_1;
input 	src0_valid;
input 	ic_fill_line_5;
output 	src_data_46;
input 	ic_fill_line_0;
input 	ic_fill_line_1;
input 	ic_fill_line_2;
input 	ic_fill_line_3;
input 	ic_fill_line_4;
input 	ic_fill_ap_offset_0;
input 	ic_fill_ap_offset_1;
input 	ic_fill_ap_offset_2;
input 	M_mem_byte_en_0;
input 	M_mem_byte_en_2;
input 	M_mem_byte_en_1;
input 	M_st_data_24;
input 	M_mem_byte_en_3;
output 	src_payload;
output 	src_data_38;
output 	src_data_41;
output 	src_data_40;
output 	src_data_39;
output 	src_data_45;
output 	src_data_44;
output 	src_data_43;
output 	src_data_42;
output 	src_payload1;
input 	M_st_data_29;
input 	M_st_data_28;
input 	M_st_data_30;
input 	M_st_data_31;
input 	M_st_data_27;
input 	M_st_data_26;
input 	M_st_data_25;
output 	src_payload2;
output 	src_data_32;
output 	src_payload3;
output 	src_payload4;
output 	src_payload5;
output 	src_data_34;
output 	src_payload6;
output 	src_data_33;
output 	src_payload7;
output 	src_data_35;
output 	src_payload8;
output 	src_payload9;
output 	src_payload10;
output 	src_payload11;
output 	src_payload12;
output 	src_payload13;
output 	src_payload14;
output 	src_payload15;
output 	src_payload16;
output 	src_payload17;
output 	src_payload18;
output 	src_payload19;
output 	src_payload20;
output 	src_payload21;
output 	src_payload22;
output 	src_payload23;
output 	src_payload24;
output 	src_payload25;
output 	src_payload26;
output 	src_payload27;
output 	src_payload28;
output 	src_payload29;
output 	src_payload30;
output 	src_payload31;
output 	src_payload32;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \arb|grant[0]~0_combout ;
wire \arb|grant[1]~1_combout ;
wire \packet_in_progress~0_combout ;
wire \packet_in_progress~q ;
wire \update_grant~0_combout ;


processor_altera_merlin_arbitrator arb(
	.reset(r_sync_rst),
	.saved_grant_0(saved_grant_0),
	.write(write),
	.src2_valid(src2_valid),
	.saved_grant_1(saved_grant_1),
	.src0_valid(src0_valid),
	.grant_0(\arb|grant[0]~0_combout ),
	.packet_in_progress(\packet_in_progress~q ),
	.grant_1(\arb|grant[1]~1_combout ),
	.clk(clk_clk));

dffeas \saved_grant[0] (
	.clk(clk_clk),
	.d(\arb|grant[0]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_grant~0_combout ),
	.q(saved_grant_0),
	.prn(vcc));
defparam \saved_grant[0] .is_wysiwyg = "true";
defparam \saved_grant[0] .power_up = "low";

dffeas \saved_grant[1] (
	.clk(clk_clk),
	.d(\arb|grant[1]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_grant~0_combout ),
	.q(saved_grant_1),
	.prn(vcc));
defparam \saved_grant[1] .is_wysiwyg = "true";
defparam \saved_grant[1] .power_up = "low";

cyclonev_lcell_comb \src_data[46] (
	.dataa(!M_alu_result_10),
	.datab(!saved_grant_0),
	.datac(!saved_grant_1),
	.datad(!ic_fill_line_5),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_46),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[46] .extended_lut = "off";
defparam \src_data[46] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[46] .shared_arith = "off";

cyclonev_lcell_comb \src_payload~0 (
	.dataa(!M_st_data_3),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~0 .extended_lut = "off";
defparam \src_payload~0 .lut_mask = 64'h7777777777777777;
defparam \src_payload~0 .shared_arith = "off";

cyclonev_lcell_comb \src_data[38] (
	.dataa(!M_alu_result_2),
	.datab(!saved_grant_0),
	.datac(!saved_grant_1),
	.datad(!ic_fill_ap_offset_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_38),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[38] .extended_lut = "off";
defparam \src_data[38] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[38] .shared_arith = "off";

cyclonev_lcell_comb \src_data[41] (
	.dataa(!M_alu_result_5),
	.datab(!saved_grant_0),
	.datac(!saved_grant_1),
	.datad(!ic_fill_line_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_41),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[41] .extended_lut = "off";
defparam \src_data[41] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[41] .shared_arith = "off";

cyclonev_lcell_comb \src_data[40] (
	.dataa(!M_alu_result_4),
	.datab(!saved_grant_0),
	.datac(!saved_grant_1),
	.datad(!ic_fill_ap_offset_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_40),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[40] .extended_lut = "off";
defparam \src_data[40] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[40] .shared_arith = "off";

cyclonev_lcell_comb \src_data[39] (
	.dataa(!M_alu_result_3),
	.datab(!saved_grant_0),
	.datac(!saved_grant_1),
	.datad(!ic_fill_ap_offset_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_39),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[39] .extended_lut = "off";
defparam \src_data[39] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[39] .shared_arith = "off";

cyclonev_lcell_comb \src_data[45] (
	.dataa(!M_alu_result_9),
	.datab(!saved_grant_0),
	.datac(!saved_grant_1),
	.datad(!ic_fill_line_4),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_45),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[45] .extended_lut = "off";
defparam \src_data[45] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[45] .shared_arith = "off";

cyclonev_lcell_comb \src_data[44] (
	.dataa(!M_alu_result_8),
	.datab(!saved_grant_0),
	.datac(!saved_grant_1),
	.datad(!ic_fill_line_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_44),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[44] .extended_lut = "off";
defparam \src_data[44] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[44] .shared_arith = "off";

cyclonev_lcell_comb \src_data[43] (
	.dataa(!M_alu_result_7),
	.datab(!saved_grant_0),
	.datac(!saved_grant_1),
	.datad(!ic_fill_line_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_43),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[43] .extended_lut = "off";
defparam \src_data[43] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[43] .shared_arith = "off";

cyclonev_lcell_comb \src_data[42] (
	.dataa(!M_alu_result_6),
	.datab(!saved_grant_0),
	.datac(!saved_grant_1),
	.datad(!ic_fill_line_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_42),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[42] .extended_lut = "off";
defparam \src_data[42] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[42] .shared_arith = "off";

cyclonev_lcell_comb \src_payload~1 (
	.dataa(!saved_grant_0),
	.datab(!hbreak_enabled),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload1),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~1 .extended_lut = "off";
defparam \src_payload~1 .lut_mask = 64'h7777777777777777;
defparam \src_payload~1 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~2 (
	.dataa(!M_st_data_0),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload2),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~2 .extended_lut = "off";
defparam \src_payload~2 .lut_mask = 64'h7777777777777777;
defparam \src_payload~2 .shared_arith = "off";

cyclonev_lcell_comb \src_data[32] (
	.dataa(!saved_grant_0),
	.datab(!saved_grant_1),
	.datac(!M_mem_byte_en_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_32),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[32] .extended_lut = "off";
defparam \src_data[32] .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \src_data[32] .shared_arith = "off";

cyclonev_lcell_comb \src_payload~3 (
	.dataa(!saved_grant_0),
	.datab(!M_st_data_16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload3),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~3 .extended_lut = "off";
defparam \src_payload~3 .lut_mask = 64'h7777777777777777;
defparam \src_payload~3 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~4 (
	.dataa(!M_st_data_1),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload4),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~4 .extended_lut = "off";
defparam \src_payload~4 .lut_mask = 64'h7777777777777777;
defparam \src_payload~4 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~5 (
	.dataa(!M_st_data_2),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload5),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~5 .extended_lut = "off";
defparam \src_payload~5 .lut_mask = 64'h7777777777777777;
defparam \src_payload~5 .shared_arith = "off";

cyclonev_lcell_comb \src_data[34] (
	.dataa(!saved_grant_0),
	.datab(!saved_grant_1),
	.datac(!M_mem_byte_en_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_34),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[34] .extended_lut = "off";
defparam \src_data[34] .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \src_data[34] .shared_arith = "off";

cyclonev_lcell_comb \src_payload~6 (
	.dataa(!M_st_data_8),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload6),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~6 .extended_lut = "off";
defparam \src_payload~6 .lut_mask = 64'h7777777777777777;
defparam \src_payload~6 .shared_arith = "off";

cyclonev_lcell_comb \src_data[33] (
	.dataa(!saved_grant_0),
	.datab(!saved_grant_1),
	.datac(!M_mem_byte_en_1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_33),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[33] .extended_lut = "off";
defparam \src_data[33] .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \src_data[33] .shared_arith = "off";

cyclonev_lcell_comb \src_payload~7 (
	.dataa(!saved_grant_0),
	.datab(!M_st_data_24),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload7),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~7 .extended_lut = "off";
defparam \src_payload~7 .lut_mask = 64'h7777777777777777;
defparam \src_payload~7 .shared_arith = "off";

cyclonev_lcell_comb \src_data[35] (
	.dataa(!saved_grant_0),
	.datab(!saved_grant_1),
	.datac(!M_mem_byte_en_3),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_35),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[35] .extended_lut = "off";
defparam \src_data[35] .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \src_data[35] .shared_arith = "off";

cyclonev_lcell_comb \src_payload~8 (
	.dataa(!saved_grant_0),
	.datab(!M_st_data_20),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload8),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~8 .extended_lut = "off";
defparam \src_payload~8 .lut_mask = 64'h7777777777777777;
defparam \src_payload~8 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~9 (
	.dataa(!saved_grant_0),
	.datab(!M_st_data_19),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload9),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~9 .extended_lut = "off";
defparam \src_payload~9 .lut_mask = 64'h7777777777777777;
defparam \src_payload~9 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~10 (
	.dataa(!M_st_data_5),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload10),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~10 .extended_lut = "off";
defparam \src_payload~10 .lut_mask = 64'h7777777777777777;
defparam \src_payload~10 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~11 (
	.dataa(!saved_grant_0),
	.datab(!M_st_data_21),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload11),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~11 .extended_lut = "off";
defparam \src_payload~11 .lut_mask = 64'h7777777777777777;
defparam \src_payload~11 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~12 (
	.dataa(!saved_grant_0),
	.datab(!M_st_data_13),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload12),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~12 .extended_lut = "off";
defparam \src_payload~12 .lut_mask = 64'h7777777777777777;
defparam \src_payload~12 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~13 (
	.dataa(!saved_grant_0),
	.datab(!M_st_data_29),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload13),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~13 .extended_lut = "off";
defparam \src_payload~13 .lut_mask = 64'h7777777777777777;
defparam \src_payload~13 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~14 (
	.dataa(!M_st_data_4),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload14),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~14 .extended_lut = "off";
defparam \src_payload~14 .lut_mask = 64'h7777777777777777;
defparam \src_payload~14 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~15 (
	.dataa(!saved_grant_0),
	.datab(!M_st_data_12),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload15),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~15 .extended_lut = "off";
defparam \src_payload~15 .lut_mask = 64'h7777777777777777;
defparam \src_payload~15 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~16 (
	.dataa(!saved_grant_0),
	.datab(!M_st_data_28),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload16),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~16 .extended_lut = "off";
defparam \src_payload~16 .lut_mask = 64'h7777777777777777;
defparam \src_payload~16 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~17 (
	.dataa(!M_st_data_6),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload17),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~17 .extended_lut = "off";
defparam \src_payload~17 .lut_mask = 64'h7777777777777777;
defparam \src_payload~17 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~18 (
	.dataa(!saved_grant_0),
	.datab(!M_st_data_22),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload18),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~18 .extended_lut = "off";
defparam \src_payload~18 .lut_mask = 64'h7777777777777777;
defparam \src_payload~18 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~19 (
	.dataa(!saved_grant_0),
	.datab(!M_st_data_14),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload19),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~19 .extended_lut = "off";
defparam \src_payload~19 .lut_mask = 64'h7777777777777777;
defparam \src_payload~19 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~20 (
	.dataa(!saved_grant_0),
	.datab(!M_st_data_30),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload20),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~20 .extended_lut = "off";
defparam \src_payload~20 .lut_mask = 64'h7777777777777777;
defparam \src_payload~20 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~21 (
	.dataa(!M_st_data_7),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload21),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~21 .extended_lut = "off";
defparam \src_payload~21 .lut_mask = 64'h7777777777777777;
defparam \src_payload~21 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~22 (
	.dataa(!saved_grant_0),
	.datab(!M_st_data_23),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload22),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~22 .extended_lut = "off";
defparam \src_payload~22 .lut_mask = 64'h7777777777777777;
defparam \src_payload~22 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~23 (
	.dataa(!saved_grant_0),
	.datab(!M_st_data_15),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload23),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~23 .extended_lut = "off";
defparam \src_payload~23 .lut_mask = 64'h7777777777777777;
defparam \src_payload~23 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~24 (
	.dataa(!saved_grant_0),
	.datab(!M_st_data_31),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload24),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~24 .extended_lut = "off";
defparam \src_payload~24 .lut_mask = 64'h7777777777777777;
defparam \src_payload~24 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~25 (
	.dataa(!saved_grant_0),
	.datab(!M_st_data_11),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload25),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~25 .extended_lut = "off";
defparam \src_payload~25 .lut_mask = 64'h7777777777777777;
defparam \src_payload~25 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~26 (
	.dataa(!saved_grant_0),
	.datab(!M_st_data_27),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload26),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~26 .extended_lut = "off";
defparam \src_payload~26 .lut_mask = 64'h7777777777777777;
defparam \src_payload~26 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~27 (
	.dataa(!saved_grant_0),
	.datab(!M_st_data_10),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload27),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~27 .extended_lut = "off";
defparam \src_payload~27 .lut_mask = 64'h7777777777777777;
defparam \src_payload~27 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~28 (
	.dataa(!saved_grant_0),
	.datab(!M_st_data_26),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload28),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~28 .extended_lut = "off";
defparam \src_payload~28 .lut_mask = 64'h7777777777777777;
defparam \src_payload~28 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~29 (
	.dataa(!saved_grant_0),
	.datab(!M_st_data_25),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload29),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~29 .extended_lut = "off";
defparam \src_payload~29 .lut_mask = 64'h7777777777777777;
defparam \src_payload~29 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~30 (
	.dataa(!M_st_data_9),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload30),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~30 .extended_lut = "off";
defparam \src_payload~30 .lut_mask = 64'h7777777777777777;
defparam \src_payload~30 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~31 (
	.dataa(!saved_grant_0),
	.datab(!M_st_data_18),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload31),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~31 .extended_lut = "off";
defparam \src_payload~31 .lut_mask = 64'h7777777777777777;
defparam \src_payload~31 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~32 (
	.dataa(!saved_grant_0),
	.datab(!M_st_data_17),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload32),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~32 .extended_lut = "off";
defparam \src_payload~32 .lut_mask = 64'h7777777777777777;
defparam \src_payload~32 .shared_arith = "off";

cyclonev_lcell_comb \packet_in_progress~0 (
	.dataa(!\update_grant~0_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\packet_in_progress~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \packet_in_progress~0 .extended_lut = "off";
defparam \packet_in_progress~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \packet_in_progress~0 .shared_arith = "off";

dffeas packet_in_progress(
	.clk(clk_clk),
	.d(\packet_in_progress~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\packet_in_progress~q ),
	.prn(vcc));
defparam packet_in_progress.is_wysiwyg = "true";
defparam packet_in_progress.power_up = "low";

cyclonev_lcell_comb \update_grant~0 (
	.dataa(!saved_grant_0),
	.datab(!write),
	.datac(!src2_valid),
	.datad(!saved_grant_1),
	.datae(!src0_valid),
	.dataf(!\packet_in_progress~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\update_grant~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \update_grant~0 .extended_lut = "off";
defparam \update_grant~0 .lut_mask = 64'hFFFFFFFF7BB7B77B;
defparam \update_grant~0 .shared_arith = "off";

endmodule

module processor_altera_merlin_arbitrator (
	reset,
	saved_grant_0,
	write,
	src2_valid,
	saved_grant_1,
	src0_valid,
	grant_0,
	packet_in_progress,
	grant_1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset;
input 	saved_grant_0;
input 	write;
input 	src2_valid;
input 	saved_grant_1;
input 	src0_valid;
output 	grant_0;
input 	packet_in_progress;
output 	grant_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \top_priority_reg[0]~1_combout ;
wire \top_priority_reg[0]~0_combout ;
wire \top_priority_reg[0]~q ;
wire \top_priority_reg[1]~q ;


cyclonev_lcell_comb \grant[0]~0 (
	.dataa(!src2_valid),
	.datab(!src0_valid),
	.datac(!\top_priority_reg[0]~q ),
	.datad(!\top_priority_reg[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(grant_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \grant[0]~0 .extended_lut = "off";
defparam \grant[0]~0 .lut_mask = 64'hFDFFFDFFFDFFFDFF;
defparam \grant[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \grant[1]~1 (
	.dataa(!src2_valid),
	.datab(!src0_valid),
	.datac(!\top_priority_reg[0]~q ),
	.datad(!\top_priority_reg[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(grant_1),
	.sumout(),
	.cout(),
	.shareout());
defparam \grant[1]~1 .extended_lut = "off";
defparam \grant[1]~1 .lut_mask = 64'hFBFFFBFFFBFFFBFF;
defparam \grant[1]~1 .shared_arith = "off";

cyclonev_lcell_comb \top_priority_reg[0]~1 (
	.dataa(!grant_1),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\top_priority_reg[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \top_priority_reg[0]~1 .extended_lut = "off";
defparam \top_priority_reg[0]~1 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \top_priority_reg[0]~1 .shared_arith = "off";

cyclonev_lcell_comb \top_priority_reg[0]~0 (
	.dataa(!saved_grant_0),
	.datab(!write),
	.datac(!src2_valid),
	.datad(!saved_grant_1),
	.datae(!src0_valid),
	.dataf(!packet_in_progress),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\top_priority_reg[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \top_priority_reg[0]~0 .extended_lut = "off";
defparam \top_priority_reg[0]~0 .lut_mask = 64'hFFFFFFFF7BB7B77B;
defparam \top_priority_reg[0]~0 .shared_arith = "off";

dffeas \top_priority_reg[0] (
	.clk(clk),
	.d(\top_priority_reg[0]~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\top_priority_reg[0]~0_combout ),
	.q(\top_priority_reg[0]~q ),
	.prn(vcc));
defparam \top_priority_reg[0] .is_wysiwyg = "true";
defparam \top_priority_reg[0] .power_up = "low";

dffeas \top_priority_reg[1] (
	.clk(clk),
	.d(grant_0),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\top_priority_reg[0]~0_combout ),
	.q(\top_priority_reg[1]~q ),
	.prn(vcc));
defparam \top_priority_reg[1] .is_wysiwyg = "true";
defparam \top_priority_reg[1] .power_up = "low";

endmodule

module processor_processor_mm_interconnect_0_cmd_mux_002_1 (
	M_st_data_8,
	M_st_data_9,
	M_st_data_16,
	M_st_data_21,
	M_st_data_13,
	M_st_data_20,
	M_st_data_12,
	M_st_data_22,
	M_st_data_14,
	M_st_data_23,
	M_st_data_15,
	M_st_data_11,
	M_st_data_10,
	M_st_data_19,
	M_st_data_18,
	M_st_data_17,
	M_st_data_0,
	r_sync_rst,
	M_alu_result_5,
	M_alu_result_4,
	M_alu_result_6,
	M_alu_result_14,
	M_alu_result_13,
	M_alu_result_12,
	M_alu_result_11,
	M_alu_result_10,
	M_alu_result_9,
	M_alu_result_8,
	M_alu_result_7,
	M_alu_result_3,
	M_alu_result_2,
	M_st_data_1,
	M_st_data_2,
	M_st_data_3,
	M_st_data_4,
	M_st_data_5,
	M_st_data_6,
	M_st_data_7,
	saved_grant_0,
	read_latency_shift_reg,
	ic_fill_tag_3,
	ic_fill_tag_2,
	ic_fill_tag_1,
	ic_fill_tag_0,
	src3_valid,
	saved_grant_1,
	src1_valid,
	ic_fill_line_5,
	ic_fill_line_0,
	ic_fill_line_1,
	ic_fill_line_2,
	ic_fill_line_3,
	ic_fill_line_4,
	src_payload,
	ic_fill_ap_offset_0,
	src_data_38,
	ic_fill_ap_offset_1,
	src_data_39,
	ic_fill_ap_offset_2,
	src_data_40,
	src_data_41,
	src_data_42,
	src_data_43,
	src_data_44,
	src_data_45,
	src_data_46,
	src_data_47,
	src_data_48,
	src_data_49,
	src_data_50,
	M_mem_byte_en_0,
	src_data_32,
	src_payload1,
	M_mem_byte_en_2,
	src_data_34,
	src_payload2,
	M_mem_byte_en_1,
	src_data_33,
	M_st_data_24,
	src_payload3,
	M_mem_byte_en_3,
	src_data_35,
	src_payload4,
	src_payload5,
	src_payload6,
	M_st_data_29,
	src_payload7,
	src_payload8,
	src_payload9,
	src_payload10,
	M_st_data_28,
	src_payload11,
	src_payload12,
	src_payload13,
	src_payload14,
	M_st_data_30,
	src_payload15,
	src_payload16,
	src_payload17,
	src_payload18,
	M_st_data_31,
	src_payload19,
	src_payload20,
	M_st_data_27,
	src_payload21,
	src_payload22,
	M_st_data_26,
	src_payload23,
	M_st_data_25,
	src_payload24,
	src_payload25,
	src_payload26,
	src_payload27,
	src_payload28,
	src_payload29,
	src_payload30,
	src_payload31,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	M_st_data_8;
input 	M_st_data_9;
input 	M_st_data_16;
input 	M_st_data_21;
input 	M_st_data_13;
input 	M_st_data_20;
input 	M_st_data_12;
input 	M_st_data_22;
input 	M_st_data_14;
input 	M_st_data_23;
input 	M_st_data_15;
input 	M_st_data_11;
input 	M_st_data_10;
input 	M_st_data_19;
input 	M_st_data_18;
input 	M_st_data_17;
input 	M_st_data_0;
input 	r_sync_rst;
input 	M_alu_result_5;
input 	M_alu_result_4;
input 	M_alu_result_6;
input 	M_alu_result_14;
input 	M_alu_result_13;
input 	M_alu_result_12;
input 	M_alu_result_11;
input 	M_alu_result_10;
input 	M_alu_result_9;
input 	M_alu_result_8;
input 	M_alu_result_7;
input 	M_alu_result_3;
input 	M_alu_result_2;
input 	M_st_data_1;
input 	M_st_data_2;
input 	M_st_data_3;
input 	M_st_data_4;
input 	M_st_data_5;
input 	M_st_data_6;
input 	M_st_data_7;
output 	saved_grant_0;
input 	read_latency_shift_reg;
input 	ic_fill_tag_3;
input 	ic_fill_tag_2;
input 	ic_fill_tag_1;
input 	ic_fill_tag_0;
input 	src3_valid;
output 	saved_grant_1;
input 	src1_valid;
input 	ic_fill_line_5;
input 	ic_fill_line_0;
input 	ic_fill_line_1;
input 	ic_fill_line_2;
input 	ic_fill_line_3;
input 	ic_fill_line_4;
output 	src_payload;
input 	ic_fill_ap_offset_0;
output 	src_data_38;
input 	ic_fill_ap_offset_1;
output 	src_data_39;
input 	ic_fill_ap_offset_2;
output 	src_data_40;
output 	src_data_41;
output 	src_data_42;
output 	src_data_43;
output 	src_data_44;
output 	src_data_45;
output 	src_data_46;
output 	src_data_47;
output 	src_data_48;
output 	src_data_49;
output 	src_data_50;
input 	M_mem_byte_en_0;
output 	src_data_32;
output 	src_payload1;
input 	M_mem_byte_en_2;
output 	src_data_34;
output 	src_payload2;
input 	M_mem_byte_en_1;
output 	src_data_33;
input 	M_st_data_24;
output 	src_payload3;
input 	M_mem_byte_en_3;
output 	src_data_35;
output 	src_payload4;
output 	src_payload5;
output 	src_payload6;
input 	M_st_data_29;
output 	src_payload7;
output 	src_payload8;
output 	src_payload9;
output 	src_payload10;
input 	M_st_data_28;
output 	src_payload11;
output 	src_payload12;
output 	src_payload13;
output 	src_payload14;
input 	M_st_data_30;
output 	src_payload15;
output 	src_payload16;
output 	src_payload17;
output 	src_payload18;
input 	M_st_data_31;
output 	src_payload19;
output 	src_payload20;
input 	M_st_data_27;
output 	src_payload21;
output 	src_payload22;
input 	M_st_data_26;
output 	src_payload23;
input 	M_st_data_25;
output 	src_payload24;
output 	src_payload25;
output 	src_payload26;
output 	src_payload27;
output 	src_payload28;
output 	src_payload29;
output 	src_payload30;
output 	src_payload31;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \arb|grant[0]~0_combout ;
wire \arb|grant[1]~1_combout ;
wire \packet_in_progress~0_combout ;
wire \packet_in_progress~q ;
wire \update_grant~0_combout ;


processor_altera_merlin_arbitrator_1 arb(
	.reset(r_sync_rst),
	.saved_grant_0(saved_grant_0),
	.read_latency_shift_reg(read_latency_shift_reg),
	.src3_valid(src3_valid),
	.saved_grant_1(saved_grant_1),
	.src1_valid(src1_valid),
	.grant_0(\arb|grant[0]~0_combout ),
	.packet_in_progress(\packet_in_progress~q ),
	.grant_1(\arb|grant[1]~1_combout ),
	.clk(clk_clk));

dffeas \saved_grant[0] (
	.clk(clk_clk),
	.d(\arb|grant[0]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_grant~0_combout ),
	.q(saved_grant_0),
	.prn(vcc));
defparam \saved_grant[0] .is_wysiwyg = "true";
defparam \saved_grant[0] .power_up = "low";

dffeas \saved_grant[1] (
	.clk(clk_clk),
	.d(\arb|grant[1]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_grant~0_combout ),
	.q(saved_grant_1),
	.prn(vcc));
defparam \saved_grant[1] .is_wysiwyg = "true";
defparam \saved_grant[1] .power_up = "low";

cyclonev_lcell_comb \src_payload~0 (
	.dataa(!M_st_data_0),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~0 .extended_lut = "off";
defparam \src_payload~0 .lut_mask = 64'h7777777777777777;
defparam \src_payload~0 .shared_arith = "off";

cyclonev_lcell_comb \src_data[38] (
	.dataa(!M_alu_result_2),
	.datab(!saved_grant_0),
	.datac(!saved_grant_1),
	.datad(!ic_fill_ap_offset_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_38),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[38] .extended_lut = "off";
defparam \src_data[38] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[38] .shared_arith = "off";

cyclonev_lcell_comb \src_data[39] (
	.dataa(!M_alu_result_3),
	.datab(!saved_grant_0),
	.datac(!saved_grant_1),
	.datad(!ic_fill_ap_offset_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_39),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[39] .extended_lut = "off";
defparam \src_data[39] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[39] .shared_arith = "off";

cyclonev_lcell_comb \src_data[40] (
	.dataa(!M_alu_result_4),
	.datab(!saved_grant_0),
	.datac(!saved_grant_1),
	.datad(!ic_fill_ap_offset_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_40),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[40] .extended_lut = "off";
defparam \src_data[40] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[40] .shared_arith = "off";

cyclonev_lcell_comb \src_data[41] (
	.dataa(!M_alu_result_5),
	.datab(!saved_grant_0),
	.datac(!saved_grant_1),
	.datad(!ic_fill_line_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_41),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[41] .extended_lut = "off";
defparam \src_data[41] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[41] .shared_arith = "off";

cyclonev_lcell_comb \src_data[42] (
	.dataa(!M_alu_result_6),
	.datab(!saved_grant_0),
	.datac(!saved_grant_1),
	.datad(!ic_fill_line_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_42),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[42] .extended_lut = "off";
defparam \src_data[42] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[42] .shared_arith = "off";

cyclonev_lcell_comb \src_data[43] (
	.dataa(!M_alu_result_7),
	.datab(!saved_grant_0),
	.datac(!saved_grant_1),
	.datad(!ic_fill_line_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_43),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[43] .extended_lut = "off";
defparam \src_data[43] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[43] .shared_arith = "off";

cyclonev_lcell_comb \src_data[44] (
	.dataa(!M_alu_result_8),
	.datab(!saved_grant_0),
	.datac(!saved_grant_1),
	.datad(!ic_fill_line_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_44),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[44] .extended_lut = "off";
defparam \src_data[44] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[44] .shared_arith = "off";

cyclonev_lcell_comb \src_data[45] (
	.dataa(!M_alu_result_9),
	.datab(!saved_grant_0),
	.datac(!saved_grant_1),
	.datad(!ic_fill_line_4),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_45),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[45] .extended_lut = "off";
defparam \src_data[45] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[45] .shared_arith = "off";

cyclonev_lcell_comb \src_data[46] (
	.dataa(!M_alu_result_10),
	.datab(!saved_grant_0),
	.datac(!saved_grant_1),
	.datad(!ic_fill_line_5),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_46),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[46] .extended_lut = "off";
defparam \src_data[46] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[46] .shared_arith = "off";

cyclonev_lcell_comb \src_data[47] (
	.dataa(!M_alu_result_11),
	.datab(!saved_grant_0),
	.datac(!ic_fill_tag_0),
	.datad(!saved_grant_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_47),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[47] .extended_lut = "off";
defparam \src_data[47] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[47] .shared_arith = "off";

cyclonev_lcell_comb \src_data[48] (
	.dataa(!M_alu_result_12),
	.datab(!saved_grant_0),
	.datac(!ic_fill_tag_1),
	.datad(!saved_grant_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_48),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[48] .extended_lut = "off";
defparam \src_data[48] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[48] .shared_arith = "off";

cyclonev_lcell_comb \src_data[49] (
	.dataa(!M_alu_result_13),
	.datab(!saved_grant_0),
	.datac(!ic_fill_tag_2),
	.datad(!saved_grant_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_49),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[49] .extended_lut = "off";
defparam \src_data[49] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[49] .shared_arith = "off";

cyclonev_lcell_comb \src_data[50] (
	.dataa(!M_alu_result_14),
	.datab(!saved_grant_0),
	.datac(!ic_fill_tag_3),
	.datad(!saved_grant_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_50),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[50] .extended_lut = "off";
defparam \src_data[50] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[50] .shared_arith = "off";

cyclonev_lcell_comb \src_data[32] (
	.dataa(!saved_grant_0),
	.datab(!saved_grant_1),
	.datac(!M_mem_byte_en_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_32),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[32] .extended_lut = "off";
defparam \src_data[32] .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \src_data[32] .shared_arith = "off";

cyclonev_lcell_comb \src_payload~1 (
	.dataa(!saved_grant_0),
	.datab(!M_st_data_16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload1),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~1 .extended_lut = "off";
defparam \src_payload~1 .lut_mask = 64'h7777777777777777;
defparam \src_payload~1 .shared_arith = "off";

cyclonev_lcell_comb \src_data[34] (
	.dataa(!saved_grant_0),
	.datab(!saved_grant_1),
	.datac(!M_mem_byte_en_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_34),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[34] .extended_lut = "off";
defparam \src_data[34] .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \src_data[34] .shared_arith = "off";

cyclonev_lcell_comb \src_payload~2 (
	.dataa(!M_st_data_8),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload2),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~2 .extended_lut = "off";
defparam \src_payload~2 .lut_mask = 64'h7777777777777777;
defparam \src_payload~2 .shared_arith = "off";

cyclonev_lcell_comb \src_data[33] (
	.dataa(!saved_grant_0),
	.datab(!saved_grant_1),
	.datac(!M_mem_byte_en_1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_33),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[33] .extended_lut = "off";
defparam \src_data[33] .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \src_data[33] .shared_arith = "off";

cyclonev_lcell_comb \src_payload~3 (
	.dataa(!saved_grant_0),
	.datab(!M_st_data_24),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload3),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~3 .extended_lut = "off";
defparam \src_payload~3 .lut_mask = 64'h7777777777777777;
defparam \src_payload~3 .shared_arith = "off";

cyclonev_lcell_comb \src_data[35] (
	.dataa(!saved_grant_0),
	.datab(!saved_grant_1),
	.datac(!M_mem_byte_en_3),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_35),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[35] .extended_lut = "off";
defparam \src_data[35] .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \src_data[35] .shared_arith = "off";

cyclonev_lcell_comb \src_payload~4 (
	.dataa(!M_st_data_5),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload4),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~4 .extended_lut = "off";
defparam \src_payload~4 .lut_mask = 64'h7777777777777777;
defparam \src_payload~4 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~5 (
	.dataa(!saved_grant_0),
	.datab(!M_st_data_21),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload5),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~5 .extended_lut = "off";
defparam \src_payload~5 .lut_mask = 64'h7777777777777777;
defparam \src_payload~5 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~6 (
	.dataa(!saved_grant_0),
	.datab(!M_st_data_13),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload6),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~6 .extended_lut = "off";
defparam \src_payload~6 .lut_mask = 64'h7777777777777777;
defparam \src_payload~6 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~7 (
	.dataa(!saved_grant_0),
	.datab(!M_st_data_29),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload7),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~7 .extended_lut = "off";
defparam \src_payload~7 .lut_mask = 64'h7777777777777777;
defparam \src_payload~7 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~8 (
	.dataa(!M_st_data_4),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload8),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~8 .extended_lut = "off";
defparam \src_payload~8 .lut_mask = 64'h7777777777777777;
defparam \src_payload~8 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~9 (
	.dataa(!saved_grant_0),
	.datab(!M_st_data_20),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload9),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~9 .extended_lut = "off";
defparam \src_payload~9 .lut_mask = 64'h7777777777777777;
defparam \src_payload~9 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~10 (
	.dataa(!saved_grant_0),
	.datab(!M_st_data_12),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload10),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~10 .extended_lut = "off";
defparam \src_payload~10 .lut_mask = 64'h7777777777777777;
defparam \src_payload~10 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~11 (
	.dataa(!saved_grant_0),
	.datab(!M_st_data_28),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload11),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~11 .extended_lut = "off";
defparam \src_payload~11 .lut_mask = 64'h7777777777777777;
defparam \src_payload~11 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~12 (
	.dataa(!M_st_data_6),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload12),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~12 .extended_lut = "off";
defparam \src_payload~12 .lut_mask = 64'h7777777777777777;
defparam \src_payload~12 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~13 (
	.dataa(!saved_grant_0),
	.datab(!M_st_data_22),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload13),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~13 .extended_lut = "off";
defparam \src_payload~13 .lut_mask = 64'h7777777777777777;
defparam \src_payload~13 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~14 (
	.dataa(!saved_grant_0),
	.datab(!M_st_data_14),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload14),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~14 .extended_lut = "off";
defparam \src_payload~14 .lut_mask = 64'h7777777777777777;
defparam \src_payload~14 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~15 (
	.dataa(!saved_grant_0),
	.datab(!M_st_data_30),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload15),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~15 .extended_lut = "off";
defparam \src_payload~15 .lut_mask = 64'h7777777777777777;
defparam \src_payload~15 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~16 (
	.dataa(!M_st_data_7),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload16),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~16 .extended_lut = "off";
defparam \src_payload~16 .lut_mask = 64'h7777777777777777;
defparam \src_payload~16 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~17 (
	.dataa(!saved_grant_0),
	.datab(!M_st_data_23),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload17),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~17 .extended_lut = "off";
defparam \src_payload~17 .lut_mask = 64'h7777777777777777;
defparam \src_payload~17 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~18 (
	.dataa(!saved_grant_0),
	.datab(!M_st_data_15),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload18),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~18 .extended_lut = "off";
defparam \src_payload~18 .lut_mask = 64'h7777777777777777;
defparam \src_payload~18 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~19 (
	.dataa(!saved_grant_0),
	.datab(!M_st_data_31),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload19),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~19 .extended_lut = "off";
defparam \src_payload~19 .lut_mask = 64'h7777777777777777;
defparam \src_payload~19 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~20 (
	.dataa(!saved_grant_0),
	.datab(!M_st_data_11),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload20),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~20 .extended_lut = "off";
defparam \src_payload~20 .lut_mask = 64'h7777777777777777;
defparam \src_payload~20 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~21 (
	.dataa(!saved_grant_0),
	.datab(!M_st_data_27),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload21),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~21 .extended_lut = "off";
defparam \src_payload~21 .lut_mask = 64'h7777777777777777;
defparam \src_payload~21 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~22 (
	.dataa(!saved_grant_0),
	.datab(!M_st_data_10),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload22),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~22 .extended_lut = "off";
defparam \src_payload~22 .lut_mask = 64'h7777777777777777;
defparam \src_payload~22 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~23 (
	.dataa(!saved_grant_0),
	.datab(!M_st_data_26),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload23),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~23 .extended_lut = "off";
defparam \src_payload~23 .lut_mask = 64'h7777777777777777;
defparam \src_payload~23 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~24 (
	.dataa(!saved_grant_0),
	.datab(!M_st_data_25),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload24),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~24 .extended_lut = "off";
defparam \src_payload~24 .lut_mask = 64'h7777777777777777;
defparam \src_payload~24 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~25 (
	.dataa(!M_st_data_9),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload25),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~25 .extended_lut = "off";
defparam \src_payload~25 .lut_mask = 64'h7777777777777777;
defparam \src_payload~25 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~26 (
	.dataa(!M_st_data_3),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload26),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~26 .extended_lut = "off";
defparam \src_payload~26 .lut_mask = 64'h7777777777777777;
defparam \src_payload~26 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~27 (
	.dataa(!saved_grant_0),
	.datab(!M_st_data_19),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload27),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~27 .extended_lut = "off";
defparam \src_payload~27 .lut_mask = 64'h7777777777777777;
defparam \src_payload~27 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~28 (
	.dataa(!M_st_data_2),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload28),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~28 .extended_lut = "off";
defparam \src_payload~28 .lut_mask = 64'h7777777777777777;
defparam \src_payload~28 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~29 (
	.dataa(!saved_grant_0),
	.datab(!M_st_data_18),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload29),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~29 .extended_lut = "off";
defparam \src_payload~29 .lut_mask = 64'h7777777777777777;
defparam \src_payload~29 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~30 (
	.dataa(!M_st_data_1),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload30),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~30 .extended_lut = "off";
defparam \src_payload~30 .lut_mask = 64'h7777777777777777;
defparam \src_payload~30 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~31 (
	.dataa(!saved_grant_0),
	.datab(!M_st_data_17),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload31),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~31 .extended_lut = "off";
defparam \src_payload~31 .lut_mask = 64'h7777777777777777;
defparam \src_payload~31 .shared_arith = "off";

cyclonev_lcell_comb \packet_in_progress~0 (
	.dataa(!\update_grant~0_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\packet_in_progress~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \packet_in_progress~0 .extended_lut = "off";
defparam \packet_in_progress~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \packet_in_progress~0 .shared_arith = "off";

dffeas packet_in_progress(
	.clk(clk_clk),
	.d(\packet_in_progress~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\packet_in_progress~q ),
	.prn(vcc));
defparam packet_in_progress.is_wysiwyg = "true";
defparam packet_in_progress.power_up = "low";

cyclonev_lcell_comb \update_grant~0 (
	.dataa(!saved_grant_0),
	.datab(!read_latency_shift_reg),
	.datac(!src3_valid),
	.datad(!saved_grant_1),
	.datae(!src1_valid),
	.dataf(!\packet_in_progress~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\update_grant~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \update_grant~0 .extended_lut = "off";
defparam \update_grant~0 .lut_mask = 64'hFFFFFFFF7BB7B77B;
defparam \update_grant~0 .shared_arith = "off";

endmodule

module processor_altera_merlin_arbitrator_1 (
	reset,
	saved_grant_0,
	read_latency_shift_reg,
	src3_valid,
	saved_grant_1,
	src1_valid,
	grant_0,
	packet_in_progress,
	grant_1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset;
input 	saved_grant_0;
input 	read_latency_shift_reg;
input 	src3_valid;
input 	saved_grant_1;
input 	src1_valid;
output 	grant_0;
input 	packet_in_progress;
output 	grant_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \top_priority_reg[0]~1_combout ;
wire \top_priority_reg[0]~0_combout ;
wire \top_priority_reg[0]~q ;
wire \top_priority_reg[1]~q ;


cyclonev_lcell_comb \grant[0]~0 (
	.dataa(!src3_valid),
	.datab(!src1_valid),
	.datac(!\top_priority_reg[0]~q ),
	.datad(!\top_priority_reg[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(grant_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \grant[0]~0 .extended_lut = "off";
defparam \grant[0]~0 .lut_mask = 64'hFDFFFDFFFDFFFDFF;
defparam \grant[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \grant[1]~1 (
	.dataa(!src3_valid),
	.datab(!src1_valid),
	.datac(!\top_priority_reg[0]~q ),
	.datad(!\top_priority_reg[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(grant_1),
	.sumout(),
	.cout(),
	.shareout());
defparam \grant[1]~1 .extended_lut = "off";
defparam \grant[1]~1 .lut_mask = 64'hFBFFFBFFFBFFFBFF;
defparam \grant[1]~1 .shared_arith = "off";

cyclonev_lcell_comb \top_priority_reg[0]~1 (
	.dataa(!grant_1),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\top_priority_reg[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \top_priority_reg[0]~1 .extended_lut = "off";
defparam \top_priority_reg[0]~1 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \top_priority_reg[0]~1 .shared_arith = "off";

cyclonev_lcell_comb \top_priority_reg[0]~0 (
	.dataa(!saved_grant_0),
	.datab(!read_latency_shift_reg),
	.datac(!src3_valid),
	.datad(!saved_grant_1),
	.datae(!src1_valid),
	.dataf(!packet_in_progress),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\top_priority_reg[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \top_priority_reg[0]~0 .extended_lut = "off";
defparam \top_priority_reg[0]~0 .lut_mask = 64'hFFFFFFFF7BB7B77B;
defparam \top_priority_reg[0]~0 .shared_arith = "off";

dffeas \top_priority_reg[0] (
	.clk(clk),
	.d(\top_priority_reg[0]~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\top_priority_reg[0]~0_combout ),
	.q(\top_priority_reg[0]~q ),
	.prn(vcc));
defparam \top_priority_reg[0] .is_wysiwyg = "true";
defparam \top_priority_reg[0] .power_up = "low";

dffeas \top_priority_reg[1] (
	.clk(clk),
	.d(grant_0),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\top_priority_reg[0]~0_combout ),
	.q(\top_priority_reg[1]~q ),
	.prn(vcc));
defparam \top_priority_reg[1] .is_wysiwyg = "true";
defparam \top_priority_reg[1] .power_up = "low";

endmodule

module processor_processor_mm_interconnect_0_router (
	M_alu_result_5,
	M_alu_result_4,
	M_alu_result_6,
	M_alu_result_16,
	M_alu_result_15,
	M_alu_result_14,
	M_alu_result_13,
	Equal1,
	M_alu_result_12,
	M_alu_result_11,
	M_alu_result_10,
	M_alu_result_9,
	M_alu_result_8,
	M_alu_result_7,
	Equal2,
	Equal4,
	M_alu_result_3,
	d_read,
	read_accepted,
	always1,
	always11,
	always12,
	Equal21,
	Equal6,
	Equal11,
	Equal61)/* synthesis synthesis_greybox=1 */;
input 	M_alu_result_5;
input 	M_alu_result_4;
input 	M_alu_result_6;
input 	M_alu_result_16;
input 	M_alu_result_15;
input 	M_alu_result_14;
input 	M_alu_result_13;
output 	Equal1;
input 	M_alu_result_12;
input 	M_alu_result_11;
input 	M_alu_result_10;
input 	M_alu_result_9;
input 	M_alu_result_8;
input 	M_alu_result_7;
output 	Equal2;
output 	Equal4;
input 	M_alu_result_3;
input 	d_read;
input 	read_accepted;
output 	always1;
output 	always11;
output 	always12;
output 	Equal21;
output 	Equal6;
output 	Equal11;
output 	Equal61;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb \Equal1~0 (
	.dataa(!M_alu_result_16),
	.datab(!M_alu_result_15),
	.datac(!M_alu_result_14),
	.datad(!M_alu_result_13),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Equal1),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal1~0 .extended_lut = "off";
defparam \Equal1~0 .lut_mask = 64'hFFFDFFFDFFFDFFFD;
defparam \Equal1~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal2~0 (
	.dataa(!M_alu_result_12),
	.datab(!M_alu_result_11),
	.datac(!M_alu_result_10),
	.datad(!M_alu_result_9),
	.datae(!M_alu_result_8),
	.dataf(!M_alu_result_7),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Equal2),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal2~0 .extended_lut = "off";
defparam \Equal2~0 .lut_mask = 64'hFFFFFFFFFFFFFFFD;
defparam \Equal2~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal4~0 (
	.dataa(!M_alu_result_5),
	.datab(!M_alu_result_4),
	.datac(!M_alu_result_6),
	.datad(!Equal1),
	.datae(!Equal2),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Equal4),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal4~0 .extended_lut = "off";
defparam \Equal4~0 .lut_mask = 64'hF7FFFFFFF7FFFFFF;
defparam \Equal4~0 .shared_arith = "off";

cyclonev_lcell_comb \always1~0 (
	.dataa(!M_alu_result_4),
	.datab(!d_read),
	.datac(!read_accepted),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(always1),
	.sumout(),
	.cout(),
	.shareout());
defparam \always1~0 .extended_lut = "off";
defparam \always1~0 .lut_mask = 64'hFBFBFBFBFBFBFBFB;
defparam \always1~0 .shared_arith = "off";

cyclonev_lcell_comb \always1~1 (
	.dataa(!M_alu_result_3),
	.datab(!M_alu_result_5),
	.datac(!M_alu_result_6),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(always11),
	.sumout(),
	.cout(),
	.shareout());
defparam \always1~1 .extended_lut = "off";
defparam \always1~1 .lut_mask = 64'hEFEFEFEFEFEFEFEF;
defparam \always1~1 .shared_arith = "off";

cyclonev_lcell_comb \always1~2 (
	.dataa(!M_alu_result_5),
	.datab(!M_alu_result_6),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(always12),
	.sumout(),
	.cout(),
	.shareout());
defparam \always1~2 .extended_lut = "off";
defparam \always1~2 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \always1~2 .shared_arith = "off";

cyclonev_lcell_comb \Equal2~1 (
	.dataa(!M_alu_result_5),
	.datab(!M_alu_result_6),
	.datac(!Equal1),
	.datad(!Equal2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Equal21),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal2~1 .extended_lut = "off";
defparam \Equal2~1 .lut_mask = 64'hEFFFEFFFEFFFEFFF;
defparam \Equal2~1 .shared_arith = "off";

cyclonev_lcell_comb \Equal6~0 (
	.dataa(!M_alu_result_3),
	.datab(!M_alu_result_5),
	.datac(!M_alu_result_4),
	.datad(!M_alu_result_6),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Equal6),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal6~0 .extended_lut = "off";
defparam \Equal6~0 .lut_mask = 64'hFDFFFDFFFDFFFDFF;
defparam \Equal6~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal1~1 (
	.dataa(!M_alu_result_12),
	.datab(!M_alu_result_11),
	.datac(!M_alu_result_16),
	.datad(!M_alu_result_15),
	.datae(!M_alu_result_14),
	.dataf(!M_alu_result_13),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Equal11),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal1~1 .extended_lut = "off";
defparam \Equal1~1 .lut_mask = 64'hFFFFFFFFFFFFFFBF;
defparam \Equal1~1 .shared_arith = "off";

cyclonev_lcell_comb \Equal6~1 (
	.dataa(!Equal1),
	.datab(!Equal2),
	.datac(!Equal6),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Equal61),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal6~1 .extended_lut = "off";
defparam \Equal6~1 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \Equal6~1 .shared_arith = "off";

endmodule

module processor_processor_mm_interconnect_0_router_001 (
	ic_fill_tag_5,
	ic_fill_tag_4,
	ic_fill_tag_3,
	ic_fill_tag_2,
	ic_fill_tag_1,
	ic_fill_tag_0,
	Equal1)/* synthesis synthesis_greybox=1 */;
input 	ic_fill_tag_5;
input 	ic_fill_tag_4;
input 	ic_fill_tag_3;
input 	ic_fill_tag_2;
input 	ic_fill_tag_1;
input 	ic_fill_tag_0;
output 	Equal1;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb \Equal1~0 (
	.dataa(!ic_fill_tag_5),
	.datab(!ic_fill_tag_4),
	.datac(!ic_fill_tag_3),
	.datad(!ic_fill_tag_2),
	.datae(!ic_fill_tag_1),
	.dataf(!ic_fill_tag_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Equal1),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal1~0 .extended_lut = "off";
defparam \Equal1~0 .lut_mask = 64'hFFFFFFFDFFFFFFFF;
defparam \Equal1~0 .shared_arith = "off";

endmodule

module processor_processor_mm_interconnect_0_rsp_demux_002 (
	read_latency_shift_reg_0,
	mem_74_0,
	mem_56_0,
	src0_valid,
	src1_valid)/* synthesis synthesis_greybox=1 */;
input 	read_latency_shift_reg_0;
input 	mem_74_0;
input 	mem_56_0;
output 	src0_valid;
output 	src1_valid;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb \src0_valid~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_74_0),
	.datac(!mem_56_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src0_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src0_valid~0 .extended_lut = "off";
defparam \src0_valid~0 .lut_mask = 64'hFDFDFDFDFDFDFDFD;
defparam \src0_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \src1_valid~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_74_0),
	.datac(!mem_56_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src1_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src1_valid~0 .extended_lut = "off";
defparam \src1_valid~0 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \src1_valid~0 .shared_arith = "off";

endmodule

module processor_processor_mm_interconnect_0_rsp_demux_002_1 (
	read_latency_shift_reg_0,
	mem_74_0,
	mem_56_0,
	src0_valid,
	src1_valid)/* synthesis synthesis_greybox=1 */;
input 	read_latency_shift_reg_0;
input 	mem_74_0;
input 	mem_56_0;
output 	src0_valid;
output 	src1_valid;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb \src0_valid~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_74_0),
	.datac(!mem_56_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src0_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src0_valid~0 .extended_lut = "off";
defparam \src0_valid~0 .lut_mask = 64'hFDFDFDFDFDFDFDFD;
defparam \src0_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \src1_valid~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_74_0),
	.datac(!mem_56_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src1_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src1_valid~0 .extended_lut = "off";
defparam \src1_valid~0 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \src1_valid~0 .shared_arith = "off";

endmodule

module processor_processor_mm_interconnect_0_rsp_mux (
	q_a_0,
	av_readdata_pre_0,
	av_readdata_pre_16,
	q_a_16,
	q_a_8,
	q_a_24,
	q_a_5,
	av_readdata_pre_5,
	q_a_21,
	av_readdata_pre_21,
	q_a_13,
	q_a_29,
	q_a_4,
	av_readdata_pre_4,
	q_a_20,
	av_readdata_pre_20,
	q_a_12,
	q_a_28,
	q_a_6,
	av_readdata_pre_6,
	q_a_22,
	av_readdata_pre_22,
	q_a_14,
	q_a_30,
	q_a_7,
	av_readdata_pre_7,
	q_a_23,
	q_a_15,
	q_a_31,
	q_a_11,
	q_a_27,
	q_a_10,
	q_a_26,
	q_a_25,
	q_a_9,
	q_a_3,
	av_readdata_pre_3,
	q_a_19,
	av_readdata_pre_19,
	q_a_2,
	av_readdata_pre_2,
	av_readdata_pre_18,
	q_a_18,
	q_a_1,
	av_readdata_pre_1,
	q_a_17,
	av_readdata_pre_17,
	read_latency_shift_reg_0,
	src0_valid,
	src0_valid1,
	read_latency_shift_reg_01,
	read_latency_shift_reg_02,
	read_latency_shift_reg_03,
	read_latency_shift_reg_04,
	WideOr11,
	av_readdata_pre_01,
	av_readdata_pre_02,
	av_readdata_pre_03,
	av_readdata_pre_30,
	av_readdata_pre_04,
	src_data_0,
	av_readdata_pre_161,
	src_payload,
	av_readdata_pre_8,
	av_readdata_pre_81,
	av_readdata_pre_82,
	av_readdata_pre_83,
	av_readdata_pre_84,
	src_data_8,
	av_readdata_pre_24,
	src_payload1,
	av_readdata_pre_51,
	av_readdata_pre_52,
	av_readdata_pre_53,
	av_readdata_pre_54,
	src_data_5,
	av_readdata_pre_211,
	src_payload2,
	av_readdata_pre_13,
	av_readdata_pre_131,
	av_readdata_pre_132,
	src_payload3,
	av_readdata_pre_29,
	src_payload4,
	av_readdata_pre_41,
	av_readdata_pre_42,
	av_readdata_pre_43,
	av_readdata_pre_44,
	src_data_4,
	av_readdata_pre_201,
	src_payload5,
	av_readdata_pre_12,
	av_readdata_pre_121,
	av_readdata_pre_122,
	src_payload6,
	av_readdata_pre_28,
	src_payload7,
	av_readdata_pre_61,
	av_readdata_pre_62,
	av_readdata_pre_63,
	av_readdata_pre_64,
	src_data_6,
	av_readdata_pre_221,
	src_payload8,
	av_readdata_pre_14,
	av_readdata_pre_141,
	av_readdata_pre_142,
	src_payload9,
	av_readdata_pre_301,
	src_payload10,
	av_readdata_pre_71,
	av_readdata_pre_72,
	av_readdata_pre_73,
	av_readdata_pre_74,
	src_data_7,
	av_readdata_pre_23,
	src_payload11,
	av_readdata_pre_15,
	av_readdata_pre_151,
	av_readdata_pre_152,
	src_payload12,
	av_readdata_pre_31,
	src_payload13,
	av_readdata_pre_11,
	av_readdata_pre_111,
	src_payload14,
	av_readdata_pre_27,
	src_payload15,
	av_readdata_pre_10,
	av_readdata_pre_101,
	av_readdata_pre_102,
	src_payload16,
	av_readdata_pre_26,
	src_payload17,
	av_readdata_pre_25,
	src_payload18,
	av_readdata_pre_9,
	av_readdata_pre_91,
	av_readdata_pre_92,
	av_readdata_pre_93,
	av_readdata_pre_94,
	src_data_9,
	av_readdata_pre_32,
	av_readdata_pre_33,
	av_readdata_pre_34,
	av_readdata_pre_35,
	src_data_3,
	av_readdata_pre_191,
	src_payload19,
	av_readdata_pre_210,
	av_readdata_pre_212,
	av_readdata_pre_213,
	av_readdata_pre_214,
	src_data_2,
	av_readdata_pre_181,
	src_payload20,
	av_readdata_pre_110,
	av_readdata_pre_112,
	av_readdata_pre_113,
	av_readdata_pre_114,
	src_data_1,
	av_readdata_pre_171,
	src_payload21)/* synthesis synthesis_greybox=1 */;
input 	q_a_0;
input 	av_readdata_pre_0;
input 	av_readdata_pre_16;
input 	q_a_16;
input 	q_a_8;
input 	q_a_24;
input 	q_a_5;
input 	av_readdata_pre_5;
input 	q_a_21;
input 	av_readdata_pre_21;
input 	q_a_13;
input 	q_a_29;
input 	q_a_4;
input 	av_readdata_pre_4;
input 	q_a_20;
input 	av_readdata_pre_20;
input 	q_a_12;
input 	q_a_28;
input 	q_a_6;
input 	av_readdata_pre_6;
input 	q_a_22;
input 	av_readdata_pre_22;
input 	q_a_14;
input 	q_a_30;
input 	q_a_7;
input 	av_readdata_pre_7;
input 	q_a_23;
input 	q_a_15;
input 	q_a_31;
input 	q_a_11;
input 	q_a_27;
input 	q_a_10;
input 	q_a_26;
input 	q_a_25;
input 	q_a_9;
input 	q_a_3;
input 	av_readdata_pre_3;
input 	q_a_19;
input 	av_readdata_pre_19;
input 	q_a_2;
input 	av_readdata_pre_2;
input 	av_readdata_pre_18;
input 	q_a_18;
input 	q_a_1;
input 	av_readdata_pre_1;
input 	q_a_17;
input 	av_readdata_pre_17;
input 	read_latency_shift_reg_0;
input 	src0_valid;
input 	src0_valid1;
input 	read_latency_shift_reg_01;
input 	read_latency_shift_reg_02;
input 	read_latency_shift_reg_03;
input 	read_latency_shift_reg_04;
output 	WideOr11;
input 	av_readdata_pre_01;
input 	av_readdata_pre_02;
input 	av_readdata_pre_03;
input 	av_readdata_pre_30;
input 	av_readdata_pre_04;
output 	src_data_0;
input 	av_readdata_pre_161;
output 	src_payload;
input 	av_readdata_pre_8;
input 	av_readdata_pre_81;
input 	av_readdata_pre_82;
input 	av_readdata_pre_83;
input 	av_readdata_pre_84;
output 	src_data_8;
input 	av_readdata_pre_24;
output 	src_payload1;
input 	av_readdata_pre_51;
input 	av_readdata_pre_52;
input 	av_readdata_pre_53;
input 	av_readdata_pre_54;
output 	src_data_5;
input 	av_readdata_pre_211;
output 	src_payload2;
input 	av_readdata_pre_13;
input 	av_readdata_pre_131;
input 	av_readdata_pre_132;
output 	src_payload3;
input 	av_readdata_pre_29;
output 	src_payload4;
input 	av_readdata_pre_41;
input 	av_readdata_pre_42;
input 	av_readdata_pre_43;
input 	av_readdata_pre_44;
output 	src_data_4;
input 	av_readdata_pre_201;
output 	src_payload5;
input 	av_readdata_pre_12;
input 	av_readdata_pre_121;
input 	av_readdata_pre_122;
output 	src_payload6;
input 	av_readdata_pre_28;
output 	src_payload7;
input 	av_readdata_pre_61;
input 	av_readdata_pre_62;
input 	av_readdata_pre_63;
input 	av_readdata_pre_64;
output 	src_data_6;
input 	av_readdata_pre_221;
output 	src_payload8;
input 	av_readdata_pre_14;
input 	av_readdata_pre_141;
input 	av_readdata_pre_142;
output 	src_payload9;
input 	av_readdata_pre_301;
output 	src_payload10;
input 	av_readdata_pre_71;
input 	av_readdata_pre_72;
input 	av_readdata_pre_73;
input 	av_readdata_pre_74;
output 	src_data_7;
input 	av_readdata_pre_23;
output 	src_payload11;
input 	av_readdata_pre_15;
input 	av_readdata_pre_151;
input 	av_readdata_pre_152;
output 	src_payload12;
input 	av_readdata_pre_31;
output 	src_payload13;
input 	av_readdata_pre_11;
input 	av_readdata_pre_111;
output 	src_payload14;
input 	av_readdata_pre_27;
output 	src_payload15;
input 	av_readdata_pre_10;
input 	av_readdata_pre_101;
input 	av_readdata_pre_102;
output 	src_payload16;
input 	av_readdata_pre_26;
output 	src_payload17;
input 	av_readdata_pre_25;
output 	src_payload18;
input 	av_readdata_pre_9;
input 	av_readdata_pre_91;
input 	av_readdata_pre_92;
input 	av_readdata_pre_93;
input 	av_readdata_pre_94;
output 	src_data_9;
input 	av_readdata_pre_32;
input 	av_readdata_pre_33;
input 	av_readdata_pre_34;
input 	av_readdata_pre_35;
output 	src_data_3;
input 	av_readdata_pre_191;
output 	src_payload19;
input 	av_readdata_pre_210;
input 	av_readdata_pre_212;
input 	av_readdata_pre_213;
input 	av_readdata_pre_214;
output 	src_data_2;
input 	av_readdata_pre_181;
output 	src_payload20;
input 	av_readdata_pre_110;
input 	av_readdata_pre_112;
input 	av_readdata_pre_113;
input 	av_readdata_pre_114;
output 	src_data_1;
input 	av_readdata_pre_171;
output 	src_payload21;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \WideOr1~0_combout ;
wire \src_payload~0_combout ;
wire \src_data[0]~0_combout ;
wire \src_data[0]~1_combout ;
wire \src_data[8]~2_combout ;
wire \src_data[8]~3_combout ;
wire \src_data[5]~4_combout ;
wire \src_data[5]~5_combout ;
wire \src_payload~3_combout ;
wire \src_payload~5_combout ;
wire \src_data[4]~6_combout ;
wire \src_data[4]~7_combout ;
wire \src_payload~8_combout ;
wire \src_payload~10_combout ;
wire \src_data[6]~8_combout ;
wire \src_data[6]~9_combout ;
wire \src_payload~13_combout ;
wire \src_payload~15_combout ;
wire \src_data[7]~10_combout ;
wire \src_data[7]~11_combout ;
wire \src_payload~19_combout ;
wire \src_payload~24_combout ;
wire \src_data[9]~12_combout ;
wire \src_data[9]~13_combout ;
wire \src_data[3]~14_combout ;
wire \src_data[3]~15_combout ;
wire \src_payload~28_combout ;
wire \src_data[2]~16_combout ;
wire \src_data[2]~17_combout ;
wire \src_data[1]~18_combout ;
wire \src_data[1]~19_combout ;
wire \src_payload~31_combout ;


cyclonev_lcell_comb WideOr1(
	.dataa(!read_latency_shift_reg_0),
	.datab(!src0_valid),
	.datac(!src0_valid1),
	.datad(!\WideOr1~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(WideOr11),
	.sumout(),
	.cout(),
	.shareout());
defparam WideOr1.extended_lut = "off";
defparam WideOr1.lut_mask = 64'hFEFFFEFFFEFFFEFF;
defparam WideOr1.shared_arith = "off";

cyclonev_lcell_comb \src_data[0] (
	.dataa(!read_latency_shift_reg_0),
	.datab(!src0_valid1),
	.datac(!q_a_0),
	.datad(!av_readdata_pre_01),
	.datae(!\src_data[0]~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[0] .extended_lut = "off";
defparam \src_data[0] .lut_mask = 64'hFFFF7FFFFFFF7FFF;
defparam \src_data[0] .shared_arith = "off";

cyclonev_lcell_comb \src_payload~1 (
	.dataa(!read_latency_shift_reg_01),
	.datab(!src0_valid),
	.datac(!src0_valid1),
	.datad(!av_readdata_pre_16),
	.datae(!av_readdata_pre_161),
	.dataf(!q_a_16),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~1 .extended_lut = "off";
defparam \src_payload~1 .lut_mask = 64'h7FFFFFFFFFFFFFFF;
defparam \src_payload~1 .shared_arith = "off";

cyclonev_lcell_comb \src_data[8] (
	.dataa(!read_latency_shift_reg_04),
	.datab(!src0_valid1),
	.datac(!q_a_8),
	.datad(!av_readdata_pre_8),
	.datae(!\src_data[8]~2_combout ),
	.dataf(!\src_data[8]~3_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_8),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[8] .extended_lut = "off";
defparam \src_data[8] .lut_mask = 64'h7FFFFFFFFFFFFFFF;
defparam \src_data[8] .shared_arith = "off";

cyclonev_lcell_comb \src_payload~2 (
	.dataa(!src0_valid),
	.datab(!src0_valid1),
	.datac(!av_readdata_pre_24),
	.datad(!q_a_24),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload1),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~2 .extended_lut = "off";
defparam \src_payload~2 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_payload~2 .shared_arith = "off";

cyclonev_lcell_comb \src_data[5] (
	.dataa(!read_latency_shift_reg_0),
	.datab(!src0_valid1),
	.datac(!q_a_5),
	.datad(!av_readdata_pre_51),
	.datae(!\src_data[5]~5_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_5),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[5] .extended_lut = "off";
defparam \src_data[5] .lut_mask = 64'hFFFF7FFFFFFF7FFF;
defparam \src_data[5] .shared_arith = "off";

cyclonev_lcell_comb \src_payload~4 (
	.dataa(!src0_valid),
	.datab(!src0_valid1),
	.datac(!av_readdata_pre_211),
	.datad(!q_a_21),
	.datae(!\src_payload~3_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload2),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~4 .extended_lut = "off";
defparam \src_payload~4 .lut_mask = 64'hFFFF7FFFFFFF7FFF;
defparam \src_payload~4 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~6 (
	.dataa(!src0_valid),
	.datab(!src0_valid1),
	.datac(!av_readdata_pre_13),
	.datad(!q_a_13),
	.datae(!\src_payload~5_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload3),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~6 .extended_lut = "off";
defparam \src_payload~6 .lut_mask = 64'hFFFF7FFFFFFF7FFF;
defparam \src_payload~6 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~7 (
	.dataa(!src0_valid),
	.datab(!src0_valid1),
	.datac(!av_readdata_pre_29),
	.datad(!q_a_29),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload4),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~7 .extended_lut = "off";
defparam \src_payload~7 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_payload~7 .shared_arith = "off";

cyclonev_lcell_comb \src_data[4] (
	.dataa(!read_latency_shift_reg_0),
	.datab(!src0_valid1),
	.datac(!q_a_4),
	.datad(!av_readdata_pre_41),
	.datae(!\src_data[4]~7_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_4),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[4] .extended_lut = "off";
defparam \src_data[4] .lut_mask = 64'hFFFF7FFFFFFF7FFF;
defparam \src_data[4] .shared_arith = "off";

cyclonev_lcell_comb \src_payload~9 (
	.dataa(!src0_valid),
	.datab(!src0_valid1),
	.datac(!av_readdata_pre_201),
	.datad(!q_a_20),
	.datae(!\src_payload~8_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload5),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~9 .extended_lut = "off";
defparam \src_payload~9 .lut_mask = 64'hFFFF7FFFFFFF7FFF;
defparam \src_payload~9 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~11 (
	.dataa(!src0_valid),
	.datab(!src0_valid1),
	.datac(!av_readdata_pre_12),
	.datad(!q_a_12),
	.datae(!\src_payload~10_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload6),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~11 .extended_lut = "off";
defparam \src_payload~11 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \src_payload~11 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~12 (
	.dataa(!src0_valid),
	.datab(!src0_valid1),
	.datac(!\src_payload~0_combout ),
	.datad(!av_readdata_pre_28),
	.datae(!q_a_28),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload7),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~12 .extended_lut = "off";
defparam \src_payload~12 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \src_payload~12 .shared_arith = "off";

cyclonev_lcell_comb \src_data[6] (
	.dataa(!read_latency_shift_reg_0),
	.datab(!src0_valid1),
	.datac(!q_a_6),
	.datad(!av_readdata_pre_61),
	.datae(!\src_data[6]~9_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_6),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[6] .extended_lut = "off";
defparam \src_data[6] .lut_mask = 64'hFFFF7FFFFFFF7FFF;
defparam \src_data[6] .shared_arith = "off";

cyclonev_lcell_comb \src_payload~14 (
	.dataa(!src0_valid),
	.datab(!src0_valid1),
	.datac(!av_readdata_pre_221),
	.datad(!q_a_22),
	.datae(!\src_payload~13_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload8),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~14 .extended_lut = "off";
defparam \src_payload~14 .lut_mask = 64'hFFFF7FFFFFFF7FFF;
defparam \src_payload~14 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~16 (
	.dataa(!src0_valid),
	.datab(!src0_valid1),
	.datac(!av_readdata_pre_14),
	.datad(!q_a_14),
	.datae(!\src_payload~15_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload9),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~16 .extended_lut = "off";
defparam \src_payload~16 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \src_payload~16 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~17 (
	.dataa(!src0_valid),
	.datab(!src0_valid1),
	.datac(!\src_payload~0_combout ),
	.datad(!av_readdata_pre_301),
	.datae(!q_a_30),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload10),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~17 .extended_lut = "off";
defparam \src_payload~17 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \src_payload~17 .shared_arith = "off";

cyclonev_lcell_comb \src_data[7] (
	.dataa(!read_latency_shift_reg_0),
	.datab(!src0_valid1),
	.datac(!q_a_7),
	.datad(!av_readdata_pre_71),
	.datae(!\src_data[7]~11_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_7),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[7] .extended_lut = "off";
defparam \src_data[7] .lut_mask = 64'hFFFF7FFFFFFF7FFF;
defparam \src_data[7] .shared_arith = "off";

cyclonev_lcell_comb \src_payload~18 (
	.dataa(!src0_valid),
	.datab(!src0_valid1),
	.datac(!av_readdata_pre_23),
	.datad(!q_a_23),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload11),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~18 .extended_lut = "off";
defparam \src_payload~18 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_payload~18 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~20 (
	.dataa(!src0_valid),
	.datab(!src0_valid1),
	.datac(!av_readdata_pre_15),
	.datad(!q_a_15),
	.datae(!\src_payload~19_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload12),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~20 .extended_lut = "off";
defparam \src_payload~20 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \src_payload~20 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~21 (
	.dataa(!src0_valid),
	.datab(!src0_valid1),
	.datac(!av_readdata_pre_31),
	.datad(!q_a_31),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload13),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~21 .extended_lut = "off";
defparam \src_payload~21 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_payload~21 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~22 (
	.dataa(!read_latency_shift_reg_03),
	.datab(!src0_valid),
	.datac(!src0_valid1),
	.datad(!av_readdata_pre_11),
	.datae(!q_a_11),
	.dataf(!av_readdata_pre_111),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload14),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~22 .extended_lut = "off";
defparam \src_payload~22 .lut_mask = 64'h7FFFFFFFFFFFFFFF;
defparam \src_payload~22 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~23 (
	.dataa(!src0_valid),
	.datab(!src0_valid1),
	.datac(!\src_payload~0_combout ),
	.datad(!av_readdata_pre_27),
	.datae(!q_a_27),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload15),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~23 .extended_lut = "off";
defparam \src_payload~23 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \src_payload~23 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~25 (
	.dataa(!src0_valid),
	.datab(!src0_valid1),
	.datac(!av_readdata_pre_10),
	.datad(!q_a_10),
	.datae(!\src_payload~24_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload16),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~25 .extended_lut = "off";
defparam \src_payload~25 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \src_payload~25 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~26 (
	.dataa(!src0_valid),
	.datab(!src0_valid1),
	.datac(!av_readdata_pre_26),
	.datad(!q_a_26),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload17),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~26 .extended_lut = "off";
defparam \src_payload~26 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_payload~26 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~27 (
	.dataa(!src0_valid),
	.datab(!src0_valid1),
	.datac(!\src_payload~0_combout ),
	.datad(!av_readdata_pre_25),
	.datae(!q_a_25),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload18),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~27 .extended_lut = "off";
defparam \src_payload~27 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \src_payload~27 .shared_arith = "off";

cyclonev_lcell_comb \src_data[9] (
	.dataa(!read_latency_shift_reg_04),
	.datab(!src0_valid1),
	.datac(!q_a_9),
	.datad(!av_readdata_pre_9),
	.datae(!\src_data[9]~12_combout ),
	.dataf(!\src_data[9]~13_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_9),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[9] .extended_lut = "off";
defparam \src_data[9] .lut_mask = 64'h7FFFFFFFFFFFFFFF;
defparam \src_data[9] .shared_arith = "off";

cyclonev_lcell_comb \src_data[3] (
	.dataa(!read_latency_shift_reg_04),
	.datab(!src0_valid1),
	.datac(!q_a_3),
	.datad(!av_readdata_pre_32),
	.datae(!\src_data[3]~14_combout ),
	.dataf(!\src_data[3]~15_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_3),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[3] .extended_lut = "off";
defparam \src_data[3] .lut_mask = 64'h7FFFFFFFFFFFFFFF;
defparam \src_data[3] .shared_arith = "off";

cyclonev_lcell_comb \src_payload~29 (
	.dataa(!src0_valid),
	.datab(!src0_valid1),
	.datac(!av_readdata_pre_191),
	.datad(!q_a_19),
	.datae(!\src_payload~28_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload19),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~29 .extended_lut = "off";
defparam \src_payload~29 .lut_mask = 64'hFFFF7FFFFFFF7FFF;
defparam \src_payload~29 .shared_arith = "off";

cyclonev_lcell_comb \src_data[2] (
	.dataa(!read_latency_shift_reg_04),
	.datab(!src0_valid1),
	.datac(!q_a_2),
	.datad(!av_readdata_pre_210),
	.datae(!\src_data[2]~16_combout ),
	.dataf(!\src_data[2]~17_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_2),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[2] .extended_lut = "off";
defparam \src_data[2] .lut_mask = 64'h7FFFFFFFFFFFFFFF;
defparam \src_data[2] .shared_arith = "off";

cyclonev_lcell_comb \src_payload~30 (
	.dataa(!read_latency_shift_reg_01),
	.datab(!src0_valid),
	.datac(!src0_valid1),
	.datad(!av_readdata_pre_18),
	.datae(!av_readdata_pre_181),
	.dataf(!q_a_18),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload20),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~30 .extended_lut = "off";
defparam \src_payload~30 .lut_mask = 64'h7FFFFFFFFFFFFFFF;
defparam \src_payload~30 .shared_arith = "off";

cyclonev_lcell_comb \src_data[1] (
	.dataa(!read_latency_shift_reg_04),
	.datab(!src0_valid1),
	.datac(!q_a_1),
	.datad(!av_readdata_pre_110),
	.datae(!\src_data[1]~18_combout ),
	.dataf(!\src_data[1]~19_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_1),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[1] .extended_lut = "off";
defparam \src_data[1] .lut_mask = 64'h7FFFFFFFFFFFFFFF;
defparam \src_data[1] .shared_arith = "off";

cyclonev_lcell_comb \src_payload~32 (
	.dataa(!src0_valid),
	.datab(!src0_valid1),
	.datac(!av_readdata_pre_171),
	.datad(!q_a_17),
	.datae(!\src_payload~31_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload21),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~32 .extended_lut = "off";
defparam \src_payload~32 .lut_mask = 64'hFFFF7FFFFFFF7FFF;
defparam \src_payload~32 .shared_arith = "off";

cyclonev_lcell_comb \WideOr1~0 (
	.dataa(!read_latency_shift_reg_01),
	.datab(!read_latency_shift_reg_02),
	.datac(!read_latency_shift_reg_03),
	.datad(!read_latency_shift_reg_04),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr1~0 .extended_lut = "off";
defparam \WideOr1~0 .lut_mask = 64'hFFFEFFFEFFFEFFFE;
defparam \WideOr1~0 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~0 (
	.dataa(!read_latency_shift_reg_02),
	.datab(!av_readdata_pre_30),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~0 .extended_lut = "off";
defparam \src_payload~0 .lut_mask = 64'h7777777777777777;
defparam \src_payload~0 .shared_arith = "off";

cyclonev_lcell_comb \src_data[0]~0 (
	.dataa(!read_latency_shift_reg_01),
	.datab(!read_latency_shift_reg_03),
	.datac(!av_readdata_pre_0),
	.datad(!\src_payload~0_combout ),
	.datae(!av_readdata_pre_04),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[0]~0 .extended_lut = "off";
defparam \src_data[0]~0 .lut_mask = 64'hFFFFFFFEFFFFFFFE;
defparam \src_data[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \src_data[0]~1 (
	.dataa(!read_latency_shift_reg_04),
	.datab(!src0_valid),
	.datac(!av_readdata_pre_02),
	.datad(!av_readdata_pre_03),
	.datae(!\src_data[0]~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[0]~1 .extended_lut = "off";
defparam \src_data[0]~1 .lut_mask = 64'hFFFEFFFFFFFEFFFF;
defparam \src_data[0]~1 .shared_arith = "off";

cyclonev_lcell_comb \src_data[8]~2 (
	.dataa(!read_latency_shift_reg_01),
	.datab(!read_latency_shift_reg_03),
	.datac(!av_readdata_pre_81),
	.datad(!av_readdata_pre_82),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[8]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[8]~2 .extended_lut = "off";
defparam \src_data[8]~2 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[8]~2 .shared_arith = "off";

cyclonev_lcell_comb \src_data[8]~3 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!src0_valid),
	.datac(!av_readdata_pre_83),
	.datad(!av_readdata_pre_84),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[8]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[8]~3 .extended_lut = "off";
defparam \src_data[8]~3 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[8]~3 .shared_arith = "off";

cyclonev_lcell_comb \src_data[5]~4 (
	.dataa(!read_latency_shift_reg_01),
	.datab(!read_latency_shift_reg_03),
	.datac(!\src_payload~0_combout ),
	.datad(!av_readdata_pre_5),
	.datae(!av_readdata_pre_54),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[5]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[5]~4 .extended_lut = "off";
defparam \src_data[5]~4 .lut_mask = 64'hFFFFFFFEFFFFFFFE;
defparam \src_data[5]~4 .shared_arith = "off";

cyclonev_lcell_comb \src_data[5]~5 (
	.dataa(!read_latency_shift_reg_04),
	.datab(!src0_valid),
	.datac(!av_readdata_pre_52),
	.datad(!av_readdata_pre_53),
	.datae(!\src_data[5]~4_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[5]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[5]~5 .extended_lut = "off";
defparam \src_data[5]~5 .lut_mask = 64'hFFFEFFFFFFFEFFFF;
defparam \src_data[5]~5 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~3 (
	.dataa(!read_latency_shift_reg_01),
	.datab(!\src_payload~0_combout ),
	.datac(!av_readdata_pre_21),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~3 .extended_lut = "off";
defparam \src_payload~3 .lut_mask = 64'hFEFEFEFEFEFEFEFE;
defparam \src_payload~3 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~5 (
	.dataa(!read_latency_shift_reg_01),
	.datab(!read_latency_shift_reg_03),
	.datac(!\src_payload~0_combout ),
	.datad(!av_readdata_pre_131),
	.datae(!av_readdata_pre_132),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~5 .extended_lut = "off";
defparam \src_payload~5 .lut_mask = 64'hFFFFFFFEFFFFFFFE;
defparam \src_payload~5 .shared_arith = "off";

cyclonev_lcell_comb \src_data[4]~6 (
	.dataa(!read_latency_shift_reg_01),
	.datab(!read_latency_shift_reg_03),
	.datac(!\src_payload~0_combout ),
	.datad(!av_readdata_pre_4),
	.datae(!av_readdata_pre_44),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[4]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[4]~6 .extended_lut = "off";
defparam \src_data[4]~6 .lut_mask = 64'hFFFFFFFEFFFFFFFE;
defparam \src_data[4]~6 .shared_arith = "off";

cyclonev_lcell_comb \src_data[4]~7 (
	.dataa(!read_latency_shift_reg_04),
	.datab(!src0_valid),
	.datac(!av_readdata_pre_42),
	.datad(!av_readdata_pre_43),
	.datae(!\src_data[4]~6_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[4]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[4]~7 .extended_lut = "off";
defparam \src_data[4]~7 .lut_mask = 64'hFFFEFFFFFFFEFFFF;
defparam \src_data[4]~7 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~8 (
	.dataa(!read_latency_shift_reg_01),
	.datab(!\src_payload~0_combout ),
	.datac(!av_readdata_pre_20),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~8 .extended_lut = "off";
defparam \src_payload~8 .lut_mask = 64'hFEFEFEFEFEFEFEFE;
defparam \src_payload~8 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~10 (
	.dataa(!read_latency_shift_reg_01),
	.datab(!read_latency_shift_reg_03),
	.datac(!av_readdata_pre_121),
	.datad(!av_readdata_pre_122),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~10 .extended_lut = "off";
defparam \src_payload~10 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_payload~10 .shared_arith = "off";

cyclonev_lcell_comb \src_data[6]~8 (
	.dataa(!read_latency_shift_reg_01),
	.datab(!read_latency_shift_reg_03),
	.datac(!\src_payload~0_combout ),
	.datad(!av_readdata_pre_6),
	.datae(!av_readdata_pre_64),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[6]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[6]~8 .extended_lut = "off";
defparam \src_data[6]~8 .lut_mask = 64'hFFFFFFFEFFFFFFFE;
defparam \src_data[6]~8 .shared_arith = "off";

cyclonev_lcell_comb \src_data[6]~9 (
	.dataa(!read_latency_shift_reg_04),
	.datab(!src0_valid),
	.datac(!av_readdata_pre_62),
	.datad(!av_readdata_pre_63),
	.datae(!\src_data[6]~8_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[6]~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[6]~9 .extended_lut = "off";
defparam \src_data[6]~9 .lut_mask = 64'hFFFEFFFFFFFEFFFF;
defparam \src_data[6]~9 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~13 (
	.dataa(!read_latency_shift_reg_01),
	.datab(!\src_payload~0_combout ),
	.datac(!av_readdata_pre_22),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~13 .extended_lut = "off";
defparam \src_payload~13 .lut_mask = 64'hFEFEFEFEFEFEFEFE;
defparam \src_payload~13 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~15 (
	.dataa(!read_latency_shift_reg_01),
	.datab(!read_latency_shift_reg_03),
	.datac(!av_readdata_pre_141),
	.datad(!av_readdata_pre_142),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~15 .extended_lut = "off";
defparam \src_payload~15 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_payload~15 .shared_arith = "off";

cyclonev_lcell_comb \src_data[7]~10 (
	.dataa(!read_latency_shift_reg_01),
	.datab(!read_latency_shift_reg_03),
	.datac(!\src_payload~0_combout ),
	.datad(!av_readdata_pre_7),
	.datae(!av_readdata_pre_74),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[7]~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[7]~10 .extended_lut = "off";
defparam \src_data[7]~10 .lut_mask = 64'hFFFFFFFEFFFFFFFE;
defparam \src_data[7]~10 .shared_arith = "off";

cyclonev_lcell_comb \src_data[7]~11 (
	.dataa(!read_latency_shift_reg_04),
	.datab(!src0_valid),
	.datac(!av_readdata_pre_72),
	.datad(!av_readdata_pre_73),
	.datae(!\src_data[7]~10_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[7]~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[7]~11 .extended_lut = "off";
defparam \src_data[7]~11 .lut_mask = 64'hFFFEFFFFFFFEFFFF;
defparam \src_data[7]~11 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~19 (
	.dataa(!read_latency_shift_reg_01),
	.datab(!read_latency_shift_reg_03),
	.datac(!av_readdata_pre_151),
	.datad(!av_readdata_pre_152),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~19 .extended_lut = "off";
defparam \src_payload~19 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_payload~19 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~24 (
	.dataa(!read_latency_shift_reg_01),
	.datab(!read_latency_shift_reg_03),
	.datac(!av_readdata_pre_101),
	.datad(!av_readdata_pre_102),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~24_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~24 .extended_lut = "off";
defparam \src_payload~24 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_payload~24 .shared_arith = "off";

cyclonev_lcell_comb \src_data[9]~12 (
	.dataa(!read_latency_shift_reg_01),
	.datab(!read_latency_shift_reg_03),
	.datac(!av_readdata_pre_91),
	.datad(!av_readdata_pre_92),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[9]~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[9]~12 .extended_lut = "off";
defparam \src_data[9]~12 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[9]~12 .shared_arith = "off";

cyclonev_lcell_comb \src_data[9]~13 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!src0_valid),
	.datac(!av_readdata_pre_93),
	.datad(!av_readdata_pre_94),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[9]~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[9]~13 .extended_lut = "off";
defparam \src_data[9]~13 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[9]~13 .shared_arith = "off";

cyclonev_lcell_comb \src_data[3]~14 (
	.dataa(!read_latency_shift_reg_01),
	.datab(!read_latency_shift_reg_03),
	.datac(!av_readdata_pre_3),
	.datad(!av_readdata_pre_33),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[3]~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[3]~14 .extended_lut = "off";
defparam \src_data[3]~14 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[3]~14 .shared_arith = "off";

cyclonev_lcell_comb \src_data[3]~15 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!src0_valid),
	.datac(!av_readdata_pre_34),
	.datad(!av_readdata_pre_35),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[3]~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[3]~15 .extended_lut = "off";
defparam \src_data[3]~15 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[3]~15 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~28 (
	.dataa(!read_latency_shift_reg_01),
	.datab(!\src_payload~0_combout ),
	.datac(!av_readdata_pre_19),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~28_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~28 .extended_lut = "off";
defparam \src_payload~28 .lut_mask = 64'hFEFEFEFEFEFEFEFE;
defparam \src_payload~28 .shared_arith = "off";

cyclonev_lcell_comb \src_data[2]~16 (
	.dataa(!read_latency_shift_reg_01),
	.datab(!read_latency_shift_reg_03),
	.datac(!av_readdata_pre_2),
	.datad(!av_readdata_pre_212),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[2]~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[2]~16 .extended_lut = "off";
defparam \src_data[2]~16 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[2]~16 .shared_arith = "off";

cyclonev_lcell_comb \src_data[2]~17 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!src0_valid),
	.datac(!av_readdata_pre_213),
	.datad(!av_readdata_pre_214),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[2]~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[2]~17 .extended_lut = "off";
defparam \src_data[2]~17 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[2]~17 .shared_arith = "off";

cyclonev_lcell_comb \src_data[1]~18 (
	.dataa(!read_latency_shift_reg_01),
	.datab(!read_latency_shift_reg_03),
	.datac(!av_readdata_pre_1),
	.datad(!av_readdata_pre_112),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[1]~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[1]~18 .extended_lut = "off";
defparam \src_data[1]~18 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[1]~18 .shared_arith = "off";

cyclonev_lcell_comb \src_data[1]~19 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!src0_valid),
	.datac(!av_readdata_pre_113),
	.datad(!av_readdata_pre_114),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_data[1]~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[1]~19 .extended_lut = "off";
defparam \src_data[1]~19 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[1]~19 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~31 (
	.dataa(!read_latency_shift_reg_01),
	.datab(!\src_payload~0_combout ),
	.datac(!av_readdata_pre_17),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~31_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~31 .extended_lut = "off";
defparam \src_payload~31 .lut_mask = 64'hFEFEFEFEFEFEFEFE;
defparam \src_payload~31 .shared_arith = "off";

endmodule

module processor_processor_mm_interconnect_0_rsp_mux_001 (
	q_a_0,
	q_a_16,
	q_a_8,
	q_a_24,
	q_a_5,
	q_a_21,
	q_a_13,
	q_a_29,
	q_a_4,
	q_a_20,
	q_a_12,
	q_a_28,
	q_a_6,
	q_a_22,
	q_a_14,
	q_a_30,
	q_a_7,
	q_a_23,
	q_a_15,
	q_a_31,
	q_a_11,
	q_a_27,
	q_a_10,
	q_a_26,
	q_a_25,
	q_a_9,
	q_a_3,
	q_a_19,
	q_a_2,
	q_a_18,
	q_a_1,
	q_a_17,
	av_readdata_pre_0,
	av_readdata_pre_16,
	av_readdata_pre_8,
	av_readdata_pre_24,
	src1_valid,
	src1_valid1,
	av_readdata_pre_5,
	av_readdata_pre_21,
	av_readdata_pre_13,
	av_readdata_pre_29,
	av_readdata_pre_4,
	av_readdata_pre_20,
	av_readdata_pre_12,
	av_readdata_pre_28,
	av_readdata_pre_6,
	av_readdata_pre_22,
	av_readdata_pre_14,
	av_readdata_pre_30,
	av_readdata_pre_7,
	av_readdata_pre_23,
	av_readdata_pre_15,
	av_readdata_pre_31,
	av_readdata_pre_11,
	av_readdata_pre_27,
	av_readdata_pre_10,
	av_readdata_pre_26,
	av_readdata_pre_25,
	av_readdata_pre_9,
	av_readdata_pre_3,
	av_readdata_pre_19,
	av_readdata_pre_2,
	av_readdata_pre_18,
	av_readdata_pre_1,
	av_readdata_pre_17,
	WideOr11,
	src_data_24,
	src_data_0,
	src_data_1,
	src_data_2,
	src_data_3,
	src_data_4,
	src_data_5,
	src_data_22,
	src_data_23,
	src_data_25,
	src_data_26,
	src_data_14,
	src_data_12,
	src_data_11,
	src_data_16,
	src_data_15,
	src_data_13,
	src_data_21,
	src_data_29,
	src_data_27,
	src_data_28,
	src_data_30,
	src_data_31,
	src_data_10,
	src_data_6,
	src_data_8,
	src_data_7,
	src_data_20,
	src_data_19,
	src_data_18,
	src_data_17,
	src_data_9)/* synthesis synthesis_greybox=1 */;
input 	q_a_0;
input 	q_a_16;
input 	q_a_8;
input 	q_a_24;
input 	q_a_5;
input 	q_a_21;
input 	q_a_13;
input 	q_a_29;
input 	q_a_4;
input 	q_a_20;
input 	q_a_12;
input 	q_a_28;
input 	q_a_6;
input 	q_a_22;
input 	q_a_14;
input 	q_a_30;
input 	q_a_7;
input 	q_a_23;
input 	q_a_15;
input 	q_a_31;
input 	q_a_11;
input 	q_a_27;
input 	q_a_10;
input 	q_a_26;
input 	q_a_25;
input 	q_a_9;
input 	q_a_3;
input 	q_a_19;
input 	q_a_2;
input 	q_a_18;
input 	q_a_1;
input 	q_a_17;
input 	av_readdata_pre_0;
input 	av_readdata_pre_16;
input 	av_readdata_pre_8;
input 	av_readdata_pre_24;
input 	src1_valid;
input 	src1_valid1;
input 	av_readdata_pre_5;
input 	av_readdata_pre_21;
input 	av_readdata_pre_13;
input 	av_readdata_pre_29;
input 	av_readdata_pre_4;
input 	av_readdata_pre_20;
input 	av_readdata_pre_12;
input 	av_readdata_pre_28;
input 	av_readdata_pre_6;
input 	av_readdata_pre_22;
input 	av_readdata_pre_14;
input 	av_readdata_pre_30;
input 	av_readdata_pre_7;
input 	av_readdata_pre_23;
input 	av_readdata_pre_15;
input 	av_readdata_pre_31;
input 	av_readdata_pre_11;
input 	av_readdata_pre_27;
input 	av_readdata_pre_10;
input 	av_readdata_pre_26;
input 	av_readdata_pre_25;
input 	av_readdata_pre_9;
input 	av_readdata_pre_3;
input 	av_readdata_pre_19;
input 	av_readdata_pre_2;
input 	av_readdata_pre_18;
input 	av_readdata_pre_1;
input 	av_readdata_pre_17;
output 	WideOr11;
output 	src_data_24;
output 	src_data_0;
output 	src_data_1;
output 	src_data_2;
output 	src_data_3;
output 	src_data_4;
output 	src_data_5;
output 	src_data_22;
output 	src_data_23;
output 	src_data_25;
output 	src_data_26;
output 	src_data_14;
output 	src_data_12;
output 	src_data_11;
output 	src_data_16;
output 	src_data_15;
output 	src_data_13;
output 	src_data_21;
output 	src_data_29;
output 	src_data_27;
output 	src_data_28;
output 	src_data_30;
output 	src_data_31;
output 	src_data_10;
output 	src_data_6;
output 	src_data_8;
output 	src_data_7;
output 	src_data_20;
output 	src_data_19;
output 	src_data_18;
output 	src_data_17;
output 	src_data_9;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb WideOr1(
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(WideOr11),
	.sumout(),
	.cout(),
	.shareout());
defparam WideOr1.extended_lut = "off";
defparam WideOr1.lut_mask = 64'h7777777777777777;
defparam WideOr1.shared_arith = "off";

cyclonev_lcell_comb \src_data[24] (
	.dataa(!av_readdata_pre_24),
	.datab(!q_a_24),
	.datac(!src1_valid),
	.datad(!src1_valid1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_24),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[24] .extended_lut = "off";
defparam \src_data[24] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[24] .shared_arith = "off";

cyclonev_lcell_comb \src_data[0] (
	.dataa(!av_readdata_pre_0),
	.datab(!q_a_0),
	.datac(!src1_valid),
	.datad(!src1_valid1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[0] .extended_lut = "off";
defparam \src_data[0] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[0] .shared_arith = "off";

cyclonev_lcell_comb \src_data[1] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!av_readdata_pre_1),
	.datad(!q_a_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_1),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[1] .extended_lut = "off";
defparam \src_data[1] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[1] .shared_arith = "off";

cyclonev_lcell_comb \src_data[2] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!av_readdata_pre_2),
	.datad(!q_a_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_2),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[2] .extended_lut = "off";
defparam \src_data[2] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[2] .shared_arith = "off";

cyclonev_lcell_comb \src_data[3] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!av_readdata_pre_3),
	.datad(!q_a_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_3),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[3] .extended_lut = "off";
defparam \src_data[3] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[3] .shared_arith = "off";

cyclonev_lcell_comb \src_data[4] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!av_readdata_pre_4),
	.datad(!q_a_4),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_4),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[4] .extended_lut = "off";
defparam \src_data[4] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[4] .shared_arith = "off";

cyclonev_lcell_comb \src_data[5] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!av_readdata_pre_5),
	.datad(!q_a_5),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_5),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[5] .extended_lut = "off";
defparam \src_data[5] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[5] .shared_arith = "off";

cyclonev_lcell_comb \src_data[22] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!av_readdata_pre_22),
	.datad(!q_a_22),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_22),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[22] .extended_lut = "off";
defparam \src_data[22] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[22] .shared_arith = "off";

cyclonev_lcell_comb \src_data[23] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!av_readdata_pre_23),
	.datad(!q_a_23),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_23),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[23] .extended_lut = "off";
defparam \src_data[23] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[23] .shared_arith = "off";

cyclonev_lcell_comb \src_data[25] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!av_readdata_pre_25),
	.datad(!q_a_25),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_25),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[25] .extended_lut = "off";
defparam \src_data[25] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[25] .shared_arith = "off";

cyclonev_lcell_comb \src_data[26] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!av_readdata_pre_26),
	.datad(!q_a_26),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_26),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[26] .extended_lut = "off";
defparam \src_data[26] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[26] .shared_arith = "off";

cyclonev_lcell_comb \src_data[14] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!av_readdata_pre_14),
	.datad(!q_a_14),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_14),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[14] .extended_lut = "off";
defparam \src_data[14] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[14] .shared_arith = "off";

cyclonev_lcell_comb \src_data[12] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!av_readdata_pre_12),
	.datad(!q_a_12),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_12),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[12] .extended_lut = "off";
defparam \src_data[12] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[12] .shared_arith = "off";

cyclonev_lcell_comb \src_data[11] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!av_readdata_pre_11),
	.datad(!q_a_11),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_11),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[11] .extended_lut = "off";
defparam \src_data[11] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[11] .shared_arith = "off";

cyclonev_lcell_comb \src_data[16] (
	.dataa(!av_readdata_pre_16),
	.datab(!q_a_16),
	.datac(!src1_valid),
	.datad(!src1_valid1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_16),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[16] .extended_lut = "off";
defparam \src_data[16] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[16] .shared_arith = "off";

cyclonev_lcell_comb \src_data[15] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!av_readdata_pre_15),
	.datad(!q_a_15),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_15),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[15] .extended_lut = "off";
defparam \src_data[15] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[15] .shared_arith = "off";

cyclonev_lcell_comb \src_data[13] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!av_readdata_pre_13),
	.datad(!q_a_13),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_13),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[13] .extended_lut = "off";
defparam \src_data[13] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[13] .shared_arith = "off";

cyclonev_lcell_comb \src_data[21] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!av_readdata_pre_21),
	.datad(!q_a_21),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_21),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[21] .extended_lut = "off";
defparam \src_data[21] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[21] .shared_arith = "off";

cyclonev_lcell_comb \src_data[29] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!av_readdata_pre_29),
	.datad(!q_a_29),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_29),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[29] .extended_lut = "off";
defparam \src_data[29] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[29] .shared_arith = "off";

cyclonev_lcell_comb \src_data[27] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!av_readdata_pre_27),
	.datad(!q_a_27),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_27),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[27] .extended_lut = "off";
defparam \src_data[27] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[27] .shared_arith = "off";

cyclonev_lcell_comb \src_data[28] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!av_readdata_pre_28),
	.datad(!q_a_28),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_28),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[28] .extended_lut = "off";
defparam \src_data[28] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[28] .shared_arith = "off";

cyclonev_lcell_comb \src_data[30] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!av_readdata_pre_30),
	.datad(!q_a_30),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_30),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[30] .extended_lut = "off";
defparam \src_data[30] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[30] .shared_arith = "off";

cyclonev_lcell_comb \src_data[31] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!av_readdata_pre_31),
	.datad(!q_a_31),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_31),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[31] .extended_lut = "off";
defparam \src_data[31] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[31] .shared_arith = "off";

cyclonev_lcell_comb \src_data[10] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!av_readdata_pre_10),
	.datad(!q_a_10),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_10),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[10] .extended_lut = "off";
defparam \src_data[10] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[10] .shared_arith = "off";

cyclonev_lcell_comb \src_data[6] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!av_readdata_pre_6),
	.datad(!q_a_6),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_6),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[6] .extended_lut = "off";
defparam \src_data[6] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[6] .shared_arith = "off";

cyclonev_lcell_comb \src_data[8] (
	.dataa(!av_readdata_pre_8),
	.datab(!q_a_8),
	.datac(!src1_valid),
	.datad(!src1_valid1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_8),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[8] .extended_lut = "off";
defparam \src_data[8] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[8] .shared_arith = "off";

cyclonev_lcell_comb \src_data[7] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!av_readdata_pre_7),
	.datad(!q_a_7),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_7),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[7] .extended_lut = "off";
defparam \src_data[7] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[7] .shared_arith = "off";

cyclonev_lcell_comb \src_data[20] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!av_readdata_pre_20),
	.datad(!q_a_20),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_20),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[20] .extended_lut = "off";
defparam \src_data[20] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[20] .shared_arith = "off";

cyclonev_lcell_comb \src_data[19] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!av_readdata_pre_19),
	.datad(!q_a_19),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_19),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[19] .extended_lut = "off";
defparam \src_data[19] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[19] .shared_arith = "off";

cyclonev_lcell_comb \src_data[18] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!av_readdata_pre_18),
	.datad(!q_a_18),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_18),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[18] .extended_lut = "off";
defparam \src_data[18] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[18] .shared_arith = "off";

cyclonev_lcell_comb \src_data[17] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!av_readdata_pre_17),
	.datad(!q_a_17),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_17),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[17] .extended_lut = "off";
defparam \src_data[17] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[17] .shared_arith = "off";

cyclonev_lcell_comb \src_data[9] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!av_readdata_pre_9),
	.datad(!q_a_9),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_9),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[9] .extended_lut = "off";
defparam \src_data[9] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[9] .shared_arith = "off";

endmodule

module processor_processor_onchip_mem (
	q_a_0,
	q_a_16,
	q_a_8,
	q_a_24,
	q_a_5,
	q_a_21,
	q_a_13,
	q_a_29,
	q_a_4,
	q_a_20,
	q_a_12,
	q_a_28,
	q_a_6,
	q_a_22,
	q_a_14,
	q_a_30,
	q_a_7,
	q_a_23,
	q_a_15,
	q_a_31,
	q_a_11,
	q_a_27,
	q_a_10,
	q_a_26,
	q_a_25,
	q_a_9,
	q_a_3,
	q_a_19,
	q_a_2,
	q_a_18,
	q_a_1,
	q_a_17,
	d_write,
	saved_grant_0,
	mem_used_1,
	src3_valid,
	saved_grant_1,
	src1_valid,
	r_early_rst,
	src_payload,
	src_data_38,
	src_data_39,
	src_data_40,
	src_data_41,
	src_data_42,
	src_data_43,
	src_data_44,
	src_data_45,
	src_data_46,
	src_data_47,
	src_data_48,
	src_data_49,
	src_data_50,
	src_data_32,
	src_payload1,
	src_data_34,
	src_payload2,
	src_data_33,
	src_payload3,
	src_data_35,
	src_payload4,
	src_payload5,
	src_payload6,
	src_payload7,
	src_payload8,
	src_payload9,
	src_payload10,
	src_payload11,
	src_payload12,
	src_payload13,
	src_payload14,
	src_payload15,
	src_payload16,
	src_payload17,
	src_payload18,
	src_payload19,
	src_payload20,
	src_payload21,
	src_payload22,
	src_payload23,
	src_payload24,
	src_payload25,
	src_payload26,
	src_payload27,
	src_payload28,
	src_payload29,
	src_payload30,
	src_payload31,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	q_a_0;
output 	q_a_16;
output 	q_a_8;
output 	q_a_24;
output 	q_a_5;
output 	q_a_21;
output 	q_a_13;
output 	q_a_29;
output 	q_a_4;
output 	q_a_20;
output 	q_a_12;
output 	q_a_28;
output 	q_a_6;
output 	q_a_22;
output 	q_a_14;
output 	q_a_30;
output 	q_a_7;
output 	q_a_23;
output 	q_a_15;
output 	q_a_31;
output 	q_a_11;
output 	q_a_27;
output 	q_a_10;
output 	q_a_26;
output 	q_a_25;
output 	q_a_9;
output 	q_a_3;
output 	q_a_19;
output 	q_a_2;
output 	q_a_18;
output 	q_a_1;
output 	q_a_17;
input 	d_write;
input 	saved_grant_0;
input 	mem_used_1;
input 	src3_valid;
input 	saved_grant_1;
input 	src1_valid;
input 	r_early_rst;
input 	src_payload;
input 	src_data_38;
input 	src_data_39;
input 	src_data_40;
input 	src_data_41;
input 	src_data_42;
input 	src_data_43;
input 	src_data_44;
input 	src_data_45;
input 	src_data_46;
input 	src_data_47;
input 	src_data_48;
input 	src_data_49;
input 	src_data_50;
input 	src_data_32;
input 	src_payload1;
input 	src_data_34;
input 	src_payload2;
input 	src_data_33;
input 	src_payload3;
input 	src_data_35;
input 	src_payload4;
input 	src_payload5;
input 	src_payload6;
input 	src_payload7;
input 	src_payload8;
input 	src_payload9;
input 	src_payload10;
input 	src_payload11;
input 	src_payload12;
input 	src_payload13;
input 	src_payload14;
input 	src_payload15;
input 	src_payload16;
input 	src_payload17;
input 	src_payload18;
input 	src_payload19;
input 	src_payload20;
input 	src_payload21;
input 	src_payload22;
input 	src_payload23;
input 	src_payload24;
input 	src_payload25;
input 	src_payload26;
input 	src_payload27;
input 	src_payload28;
input 	src_payload29;
input 	src_payload30;
input 	src_payload31;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \wren~0_combout ;


processor_altsyncram_6 the_altsyncram(
	.q_a({q_a_31,q_a_30,q_a_29,q_a_28,q_a_27,q_a_26,q_a_25,q_a_24,q_a_23,q_a_22,q_a_21,q_a_20,q_a_19,q_a_18,q_a_17,q_a_16,q_a_15,q_a_14,q_a_13,q_a_12,q_a_11,q_a_10,q_a_9,q_a_8,q_a_7,q_a_6,q_a_5,q_a_4,q_a_3,q_a_2,q_a_1,q_a_0}),
	.clocken0(r_early_rst),
	.wren_a(\wren~0_combout ),
	.data_a({src_payload19,src_payload15,src_payload7,src_payload11,src_payload21,src_payload23,src_payload24,src_payload3,src_payload17,src_payload13,src_payload5,src_payload9,src_payload27,src_payload29,src_payload31,src_payload1,src_payload18,src_payload14,src_payload6,src_payload10,
src_payload20,src_payload22,src_payload25,src_payload2,src_payload16,src_payload12,src_payload4,src_payload8,src_payload26,src_payload28,src_payload30,src_payload}),
	.address_a({src_data_50,src_data_49,src_data_48,src_data_47,src_data_46,src_data_45,src_data_44,src_data_43,src_data_42,src_data_41,src_data_40,src_data_39,src_data_38}),
	.byteena_a({src_data_35,src_data_34,src_data_33,src_data_32}),
	.clock0(clk_clk));

cyclonev_lcell_comb \wren~0 (
	.dataa(!d_write),
	.datab(!saved_grant_0),
	.datac(!mem_used_1),
	.datad(!src3_valid),
	.datae(!saved_grant_1),
	.dataf(!src1_valid),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wren~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wren~0 .extended_lut = "off";
defparam \wren~0 .lut_mask = 64'hFFFFFFFFFFFFFFEF;
defparam \wren~0 .shared_arith = "off";

endmodule

module processor_altsyncram_6 (
	q_a,
	clocken0,
	wren_a,
	data_a,
	address_a,
	byteena_a,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[31:0] q_a;
input 	clocken0;
input 	wren_a;
input 	[31:0] data_a;
input 	[12:0] address_a;
input 	[3:0] byteena_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



processor_altsyncram_02n1 auto_generated(
	.q_a({q_a[31],q_a[30],q_a[29],q_a[28],q_a[27],q_a[26],q_a[25],q_a[24],q_a[23],q_a[22],q_a[21],q_a[20],q_a[19],q_a[18],q_a[17],q_a[16],q_a[15],q_a[14],q_a[13],q_a[12],q_a[11],q_a[10],q_a[9],q_a[8],q_a[7],q_a[6],q_a[5],q_a[4],q_a[3],q_a[2],q_a[1],q_a[0]}),
	.clocken0(clocken0),
	.wren_a(wren_a),
	.data_a({data_a[31],data_a[30],data_a[29],data_a[28],data_a[27],data_a[26],data_a[25],data_a[24],data_a[23],data_a[22],data_a[21],data_a[20],data_a[19],data_a[18],data_a[17],data_a[16],data_a[15],data_a[14],data_a[13],data_a[12],data_a[11],data_a[10],data_a[9],data_a[8],data_a[7],data_a[6],data_a[5],data_a[4],data_a[3],data_a[2],data_a[1],data_a[0]}),
	.address_a({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.byteena_a({byteena_a[3],byteena_a[2],byteena_a[1],byteena_a[0]}),
	.clock0(clock0));

endmodule

module processor_altsyncram_02n1 (
	q_a,
	clocken0,
	wren_a,
	data_a,
	address_a,
	byteena_a,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[31:0] q_a;
input 	clocken0;
input 	wren_a;
input 	[31:0] data_a;
input 	[12:0] address_a;
input 	[3:0] byteena_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a0_PORTADATAOUT_bus;
wire [143:0] ram_block1a16_PORTADATAOUT_bus;
wire [143:0] ram_block1a8_PORTADATAOUT_bus;
wire [143:0] ram_block1a24_PORTADATAOUT_bus;
wire [143:0] ram_block1a5_PORTADATAOUT_bus;
wire [143:0] ram_block1a21_PORTADATAOUT_bus;
wire [143:0] ram_block1a13_PORTADATAOUT_bus;
wire [143:0] ram_block1a29_PORTADATAOUT_bus;
wire [143:0] ram_block1a4_PORTADATAOUT_bus;
wire [143:0] ram_block1a20_PORTADATAOUT_bus;
wire [143:0] ram_block1a12_PORTADATAOUT_bus;
wire [143:0] ram_block1a28_PORTADATAOUT_bus;
wire [143:0] ram_block1a6_PORTADATAOUT_bus;
wire [143:0] ram_block1a22_PORTADATAOUT_bus;
wire [143:0] ram_block1a14_PORTADATAOUT_bus;
wire [143:0] ram_block1a30_PORTADATAOUT_bus;
wire [143:0] ram_block1a7_PORTADATAOUT_bus;
wire [143:0] ram_block1a23_PORTADATAOUT_bus;
wire [143:0] ram_block1a15_PORTADATAOUT_bus;
wire [143:0] ram_block1a31_PORTADATAOUT_bus;
wire [143:0] ram_block1a11_PORTADATAOUT_bus;
wire [143:0] ram_block1a27_PORTADATAOUT_bus;
wire [143:0] ram_block1a10_PORTADATAOUT_bus;
wire [143:0] ram_block1a26_PORTADATAOUT_bus;
wire [143:0] ram_block1a25_PORTADATAOUT_bus;
wire [143:0] ram_block1a9_PORTADATAOUT_bus;
wire [143:0] ram_block1a3_PORTADATAOUT_bus;
wire [143:0] ram_block1a19_PORTADATAOUT_bus;
wire [143:0] ram_block1a2_PORTADATAOUT_bus;
wire [143:0] ram_block1a18_PORTADATAOUT_bus;
wire [143:0] ram_block1a1_PORTADATAOUT_bus;
wire [143:0] ram_block1a17_PORTADATAOUT_bus;

assign q_a[0] = ram_block1a0_PORTADATAOUT_bus[0];

assign q_a[16] = ram_block1a16_PORTADATAOUT_bus[0];

assign q_a[8] = ram_block1a8_PORTADATAOUT_bus[0];

assign q_a[24] = ram_block1a24_PORTADATAOUT_bus[0];

assign q_a[5] = ram_block1a5_PORTADATAOUT_bus[0];

assign q_a[21] = ram_block1a21_PORTADATAOUT_bus[0];

assign q_a[13] = ram_block1a13_PORTADATAOUT_bus[0];

assign q_a[29] = ram_block1a29_PORTADATAOUT_bus[0];

assign q_a[4] = ram_block1a4_PORTADATAOUT_bus[0];

assign q_a[20] = ram_block1a20_PORTADATAOUT_bus[0];

assign q_a[12] = ram_block1a12_PORTADATAOUT_bus[0];

assign q_a[28] = ram_block1a28_PORTADATAOUT_bus[0];

assign q_a[6] = ram_block1a6_PORTADATAOUT_bus[0];

assign q_a[22] = ram_block1a22_PORTADATAOUT_bus[0];

assign q_a[14] = ram_block1a14_PORTADATAOUT_bus[0];

assign q_a[30] = ram_block1a30_PORTADATAOUT_bus[0];

assign q_a[7] = ram_block1a7_PORTADATAOUT_bus[0];

assign q_a[23] = ram_block1a23_PORTADATAOUT_bus[0];

assign q_a[15] = ram_block1a15_PORTADATAOUT_bus[0];

assign q_a[31] = ram_block1a31_PORTADATAOUT_bus[0];

assign q_a[11] = ram_block1a11_PORTADATAOUT_bus[0];

assign q_a[27] = ram_block1a27_PORTADATAOUT_bus[0];

assign q_a[10] = ram_block1a10_PORTADATAOUT_bus[0];

assign q_a[26] = ram_block1a26_PORTADATAOUT_bus[0];

assign q_a[25] = ram_block1a25_PORTADATAOUT_bus[0];

assign q_a[9] = ram_block1a9_PORTADATAOUT_bus[0];

assign q_a[3] = ram_block1a3_PORTADATAOUT_bus[0];

assign q_a[19] = ram_block1a19_PORTADATAOUT_bus[0];

assign q_a[2] = ram_block1a2_PORTADATAOUT_bus[0];

assign q_a[18] = ram_block1a18_PORTADATAOUT_bus[0];

assign q_a[1] = ram_block1a1_PORTADATAOUT_bus[0];

assign q_a[17] = ram_block1a17_PORTADATAOUT_bus[0];

cyclonev_ram_block ram_block1a0(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a0_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.clk0_input_clock_enable = "ena0";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.init_file = "processor_onchip_mem.hex";
defparam ram_block1a0.init_file_layout = "port_a";
defparam ram_block1a0.logical_ram_name = "processor_onchip_mem:onchip_mem|altsyncram:the_altsyncram|altsyncram_02n1:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.operation_mode = "single_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 13;
defparam ram_block1a0.port_a_byte_enable_mask_width = 1;
defparam ram_block1a0.port_a_byte_size = 1;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 5119;
defparam ram_block1a0.port_a_logical_ram_depth = 5120;
defparam ram_block1a0.port_a_logical_ram_width = 32;
defparam ram_block1a0.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a0.ram_block_type = "auto";
defparam ram_block1a0.mem_init2 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a0.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a0.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a16(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a16_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a16.clk0_core_clock_enable = "ena0";
defparam ram_block1a16.clk0_input_clock_enable = "ena0";
defparam ram_block1a16.data_interleave_offset_in_bits = 1;
defparam ram_block1a16.data_interleave_width_in_bits = 1;
defparam ram_block1a16.init_file = "processor_onchip_mem.hex";
defparam ram_block1a16.init_file_layout = "port_a";
defparam ram_block1a16.logical_ram_name = "processor_onchip_mem:onchip_mem|altsyncram:the_altsyncram|altsyncram_02n1:auto_generated|ALTSYNCRAM";
defparam ram_block1a16.operation_mode = "single_port";
defparam ram_block1a16.port_a_address_clear = "none";
defparam ram_block1a16.port_a_address_width = 13;
defparam ram_block1a16.port_a_byte_enable_mask_width = 1;
defparam ram_block1a16.port_a_byte_size = 1;
defparam ram_block1a16.port_a_data_out_clear = "none";
defparam ram_block1a16.port_a_data_out_clock = "none";
defparam ram_block1a16.port_a_data_width = 1;
defparam ram_block1a16.port_a_first_address = 0;
defparam ram_block1a16.port_a_first_bit_number = 16;
defparam ram_block1a16.port_a_last_address = 5119;
defparam ram_block1a16.port_a_logical_ram_depth = 5120;
defparam ram_block1a16.port_a_logical_ram_width = 32;
defparam ram_block1a16.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a16.ram_block_type = "auto";
defparam ram_block1a16.mem_init2 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a16.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a16.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a8(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a8_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a8.clk0_core_clock_enable = "ena0";
defparam ram_block1a8.clk0_input_clock_enable = "ena0";
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.init_file = "processor_onchip_mem.hex";
defparam ram_block1a8.init_file_layout = "port_a";
defparam ram_block1a8.logical_ram_name = "processor_onchip_mem:onchip_mem|altsyncram:the_altsyncram|altsyncram_02n1:auto_generated|ALTSYNCRAM";
defparam ram_block1a8.operation_mode = "single_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 13;
defparam ram_block1a8.port_a_byte_enable_mask_width = 1;
defparam ram_block1a8.port_a_byte_size = 1;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 5119;
defparam ram_block1a8.port_a_logical_ram_depth = 5120;
defparam ram_block1a8.port_a_logical_ram_width = 32;
defparam ram_block1a8.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a8.ram_block_type = "auto";
defparam ram_block1a8.mem_init2 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a8.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a8.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a24(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[24]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a24_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a24.clk0_core_clock_enable = "ena0";
defparam ram_block1a24.clk0_input_clock_enable = "ena0";
defparam ram_block1a24.data_interleave_offset_in_bits = 1;
defparam ram_block1a24.data_interleave_width_in_bits = 1;
defparam ram_block1a24.init_file = "processor_onchip_mem.hex";
defparam ram_block1a24.init_file_layout = "port_a";
defparam ram_block1a24.logical_ram_name = "processor_onchip_mem:onchip_mem|altsyncram:the_altsyncram|altsyncram_02n1:auto_generated|ALTSYNCRAM";
defparam ram_block1a24.operation_mode = "single_port";
defparam ram_block1a24.port_a_address_clear = "none";
defparam ram_block1a24.port_a_address_width = 13;
defparam ram_block1a24.port_a_byte_enable_mask_width = 1;
defparam ram_block1a24.port_a_byte_size = 1;
defparam ram_block1a24.port_a_data_out_clear = "none";
defparam ram_block1a24.port_a_data_out_clock = "none";
defparam ram_block1a24.port_a_data_width = 1;
defparam ram_block1a24.port_a_first_address = 0;
defparam ram_block1a24.port_a_first_bit_number = 24;
defparam ram_block1a24.port_a_last_address = 5119;
defparam ram_block1a24.port_a_logical_ram_depth = 5120;
defparam ram_block1a24.port_a_logical_ram_width = 32;
defparam ram_block1a24.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a24.ram_block_type = "auto";
defparam ram_block1a24.mem_init2 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a24.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a24.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a5(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a5_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a5.clk0_core_clock_enable = "ena0";
defparam ram_block1a5.clk0_input_clock_enable = "ena0";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.init_file = "processor_onchip_mem.hex";
defparam ram_block1a5.init_file_layout = "port_a";
defparam ram_block1a5.logical_ram_name = "processor_onchip_mem:onchip_mem|altsyncram:the_altsyncram|altsyncram_02n1:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.operation_mode = "single_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 13;
defparam ram_block1a5.port_a_byte_enable_mask_width = 1;
defparam ram_block1a5.port_a_byte_size = 1;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 5119;
defparam ram_block1a5.port_a_logical_ram_depth = 5120;
defparam ram_block1a5.port_a_logical_ram_width = 32;
defparam ram_block1a5.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a5.ram_block_type = "auto";
defparam ram_block1a5.mem_init2 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a5.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a5.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a21(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[21]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a21_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a21.clk0_core_clock_enable = "ena0";
defparam ram_block1a21.clk0_input_clock_enable = "ena0";
defparam ram_block1a21.data_interleave_offset_in_bits = 1;
defparam ram_block1a21.data_interleave_width_in_bits = 1;
defparam ram_block1a21.init_file = "processor_onchip_mem.hex";
defparam ram_block1a21.init_file_layout = "port_a";
defparam ram_block1a21.logical_ram_name = "processor_onchip_mem:onchip_mem|altsyncram:the_altsyncram|altsyncram_02n1:auto_generated|ALTSYNCRAM";
defparam ram_block1a21.operation_mode = "single_port";
defparam ram_block1a21.port_a_address_clear = "none";
defparam ram_block1a21.port_a_address_width = 13;
defparam ram_block1a21.port_a_byte_enable_mask_width = 1;
defparam ram_block1a21.port_a_byte_size = 1;
defparam ram_block1a21.port_a_data_out_clear = "none";
defparam ram_block1a21.port_a_data_out_clock = "none";
defparam ram_block1a21.port_a_data_width = 1;
defparam ram_block1a21.port_a_first_address = 0;
defparam ram_block1a21.port_a_first_bit_number = 21;
defparam ram_block1a21.port_a_last_address = 5119;
defparam ram_block1a21.port_a_logical_ram_depth = 5120;
defparam ram_block1a21.port_a_logical_ram_width = 32;
defparam ram_block1a21.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a21.ram_block_type = "auto";
defparam ram_block1a21.mem_init2 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a21.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a21.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a13(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a13_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a13.clk0_core_clock_enable = "ena0";
defparam ram_block1a13.clk0_input_clock_enable = "ena0";
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.init_file = "processor_onchip_mem.hex";
defparam ram_block1a13.init_file_layout = "port_a";
defparam ram_block1a13.logical_ram_name = "processor_onchip_mem:onchip_mem|altsyncram:the_altsyncram|altsyncram_02n1:auto_generated|ALTSYNCRAM";
defparam ram_block1a13.operation_mode = "single_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 13;
defparam ram_block1a13.port_a_byte_enable_mask_width = 1;
defparam ram_block1a13.port_a_byte_size = 1;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 5119;
defparam ram_block1a13.port_a_logical_ram_depth = 5120;
defparam ram_block1a13.port_a_logical_ram_width = 32;
defparam ram_block1a13.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a13.ram_block_type = "auto";
defparam ram_block1a13.mem_init2 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a13.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a13.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a29(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[29]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a29_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a29.clk0_core_clock_enable = "ena0";
defparam ram_block1a29.clk0_input_clock_enable = "ena0";
defparam ram_block1a29.data_interleave_offset_in_bits = 1;
defparam ram_block1a29.data_interleave_width_in_bits = 1;
defparam ram_block1a29.init_file = "processor_onchip_mem.hex";
defparam ram_block1a29.init_file_layout = "port_a";
defparam ram_block1a29.logical_ram_name = "processor_onchip_mem:onchip_mem|altsyncram:the_altsyncram|altsyncram_02n1:auto_generated|ALTSYNCRAM";
defparam ram_block1a29.operation_mode = "single_port";
defparam ram_block1a29.port_a_address_clear = "none";
defparam ram_block1a29.port_a_address_width = 13;
defparam ram_block1a29.port_a_byte_enable_mask_width = 1;
defparam ram_block1a29.port_a_byte_size = 1;
defparam ram_block1a29.port_a_data_out_clear = "none";
defparam ram_block1a29.port_a_data_out_clock = "none";
defparam ram_block1a29.port_a_data_width = 1;
defparam ram_block1a29.port_a_first_address = 0;
defparam ram_block1a29.port_a_first_bit_number = 29;
defparam ram_block1a29.port_a_last_address = 5119;
defparam ram_block1a29.port_a_logical_ram_depth = 5120;
defparam ram_block1a29.port_a_logical_ram_width = 32;
defparam ram_block1a29.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a29.ram_block_type = "auto";
defparam ram_block1a29.mem_init2 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a29.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a29.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a4(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a4_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a4.clk0_core_clock_enable = "ena0";
defparam ram_block1a4.clk0_input_clock_enable = "ena0";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.init_file = "processor_onchip_mem.hex";
defparam ram_block1a4.init_file_layout = "port_a";
defparam ram_block1a4.logical_ram_name = "processor_onchip_mem:onchip_mem|altsyncram:the_altsyncram|altsyncram_02n1:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.operation_mode = "single_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 13;
defparam ram_block1a4.port_a_byte_enable_mask_width = 1;
defparam ram_block1a4.port_a_byte_size = 1;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 5119;
defparam ram_block1a4.port_a_logical_ram_depth = 5120;
defparam ram_block1a4.port_a_logical_ram_width = 32;
defparam ram_block1a4.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a4.ram_block_type = "auto";
defparam ram_block1a4.mem_init2 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a4.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a4.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a20(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[20]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a20_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a20.clk0_core_clock_enable = "ena0";
defparam ram_block1a20.clk0_input_clock_enable = "ena0";
defparam ram_block1a20.data_interleave_offset_in_bits = 1;
defparam ram_block1a20.data_interleave_width_in_bits = 1;
defparam ram_block1a20.init_file = "processor_onchip_mem.hex";
defparam ram_block1a20.init_file_layout = "port_a";
defparam ram_block1a20.logical_ram_name = "processor_onchip_mem:onchip_mem|altsyncram:the_altsyncram|altsyncram_02n1:auto_generated|ALTSYNCRAM";
defparam ram_block1a20.operation_mode = "single_port";
defparam ram_block1a20.port_a_address_clear = "none";
defparam ram_block1a20.port_a_address_width = 13;
defparam ram_block1a20.port_a_byte_enable_mask_width = 1;
defparam ram_block1a20.port_a_byte_size = 1;
defparam ram_block1a20.port_a_data_out_clear = "none";
defparam ram_block1a20.port_a_data_out_clock = "none";
defparam ram_block1a20.port_a_data_width = 1;
defparam ram_block1a20.port_a_first_address = 0;
defparam ram_block1a20.port_a_first_bit_number = 20;
defparam ram_block1a20.port_a_last_address = 5119;
defparam ram_block1a20.port_a_logical_ram_depth = 5120;
defparam ram_block1a20.port_a_logical_ram_width = 32;
defparam ram_block1a20.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a20.ram_block_type = "auto";
defparam ram_block1a20.mem_init2 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a20.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a20.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a12(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a12_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a12.clk0_core_clock_enable = "ena0";
defparam ram_block1a12.clk0_input_clock_enable = "ena0";
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.init_file = "processor_onchip_mem.hex";
defparam ram_block1a12.init_file_layout = "port_a";
defparam ram_block1a12.logical_ram_name = "processor_onchip_mem:onchip_mem|altsyncram:the_altsyncram|altsyncram_02n1:auto_generated|ALTSYNCRAM";
defparam ram_block1a12.operation_mode = "single_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 13;
defparam ram_block1a12.port_a_byte_enable_mask_width = 1;
defparam ram_block1a12.port_a_byte_size = 1;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 5119;
defparam ram_block1a12.port_a_logical_ram_depth = 5120;
defparam ram_block1a12.port_a_logical_ram_width = 32;
defparam ram_block1a12.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a12.ram_block_type = "auto";
defparam ram_block1a12.mem_init2 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a12.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a12.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a28(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[28]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a28_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a28.clk0_core_clock_enable = "ena0";
defparam ram_block1a28.clk0_input_clock_enable = "ena0";
defparam ram_block1a28.data_interleave_offset_in_bits = 1;
defparam ram_block1a28.data_interleave_width_in_bits = 1;
defparam ram_block1a28.init_file = "processor_onchip_mem.hex";
defparam ram_block1a28.init_file_layout = "port_a";
defparam ram_block1a28.logical_ram_name = "processor_onchip_mem:onchip_mem|altsyncram:the_altsyncram|altsyncram_02n1:auto_generated|ALTSYNCRAM";
defparam ram_block1a28.operation_mode = "single_port";
defparam ram_block1a28.port_a_address_clear = "none";
defparam ram_block1a28.port_a_address_width = 13;
defparam ram_block1a28.port_a_byte_enable_mask_width = 1;
defparam ram_block1a28.port_a_byte_size = 1;
defparam ram_block1a28.port_a_data_out_clear = "none";
defparam ram_block1a28.port_a_data_out_clock = "none";
defparam ram_block1a28.port_a_data_width = 1;
defparam ram_block1a28.port_a_first_address = 0;
defparam ram_block1a28.port_a_first_bit_number = 28;
defparam ram_block1a28.port_a_last_address = 5119;
defparam ram_block1a28.port_a_logical_ram_depth = 5120;
defparam ram_block1a28.port_a_logical_ram_width = 32;
defparam ram_block1a28.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a28.ram_block_type = "auto";
defparam ram_block1a28.mem_init2 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a28.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a28.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a6(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a6_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a6.clk0_core_clock_enable = "ena0";
defparam ram_block1a6.clk0_input_clock_enable = "ena0";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.init_file = "processor_onchip_mem.hex";
defparam ram_block1a6.init_file_layout = "port_a";
defparam ram_block1a6.logical_ram_name = "processor_onchip_mem:onchip_mem|altsyncram:the_altsyncram|altsyncram_02n1:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.operation_mode = "single_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 13;
defparam ram_block1a6.port_a_byte_enable_mask_width = 1;
defparam ram_block1a6.port_a_byte_size = 1;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 5119;
defparam ram_block1a6.port_a_logical_ram_depth = 5120;
defparam ram_block1a6.port_a_logical_ram_width = 32;
defparam ram_block1a6.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a6.ram_block_type = "auto";
defparam ram_block1a6.mem_init2 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a6.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a6.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a22(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[22]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a22_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a22.clk0_core_clock_enable = "ena0";
defparam ram_block1a22.clk0_input_clock_enable = "ena0";
defparam ram_block1a22.data_interleave_offset_in_bits = 1;
defparam ram_block1a22.data_interleave_width_in_bits = 1;
defparam ram_block1a22.init_file = "processor_onchip_mem.hex";
defparam ram_block1a22.init_file_layout = "port_a";
defparam ram_block1a22.logical_ram_name = "processor_onchip_mem:onchip_mem|altsyncram:the_altsyncram|altsyncram_02n1:auto_generated|ALTSYNCRAM";
defparam ram_block1a22.operation_mode = "single_port";
defparam ram_block1a22.port_a_address_clear = "none";
defparam ram_block1a22.port_a_address_width = 13;
defparam ram_block1a22.port_a_byte_enable_mask_width = 1;
defparam ram_block1a22.port_a_byte_size = 1;
defparam ram_block1a22.port_a_data_out_clear = "none";
defparam ram_block1a22.port_a_data_out_clock = "none";
defparam ram_block1a22.port_a_data_width = 1;
defparam ram_block1a22.port_a_first_address = 0;
defparam ram_block1a22.port_a_first_bit_number = 22;
defparam ram_block1a22.port_a_last_address = 5119;
defparam ram_block1a22.port_a_logical_ram_depth = 5120;
defparam ram_block1a22.port_a_logical_ram_width = 32;
defparam ram_block1a22.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a22.ram_block_type = "auto";
defparam ram_block1a22.mem_init2 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a22.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a22.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a14(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a14_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a14.clk0_core_clock_enable = "ena0";
defparam ram_block1a14.clk0_input_clock_enable = "ena0";
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.init_file = "processor_onchip_mem.hex";
defparam ram_block1a14.init_file_layout = "port_a";
defparam ram_block1a14.logical_ram_name = "processor_onchip_mem:onchip_mem|altsyncram:the_altsyncram|altsyncram_02n1:auto_generated|ALTSYNCRAM";
defparam ram_block1a14.operation_mode = "single_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 13;
defparam ram_block1a14.port_a_byte_enable_mask_width = 1;
defparam ram_block1a14.port_a_byte_size = 1;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 5119;
defparam ram_block1a14.port_a_logical_ram_depth = 5120;
defparam ram_block1a14.port_a_logical_ram_width = 32;
defparam ram_block1a14.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a14.ram_block_type = "auto";
defparam ram_block1a14.mem_init2 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a14.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a14.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a30(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[30]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a30_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a30.clk0_core_clock_enable = "ena0";
defparam ram_block1a30.clk0_input_clock_enable = "ena0";
defparam ram_block1a30.data_interleave_offset_in_bits = 1;
defparam ram_block1a30.data_interleave_width_in_bits = 1;
defparam ram_block1a30.init_file = "processor_onchip_mem.hex";
defparam ram_block1a30.init_file_layout = "port_a";
defparam ram_block1a30.logical_ram_name = "processor_onchip_mem:onchip_mem|altsyncram:the_altsyncram|altsyncram_02n1:auto_generated|ALTSYNCRAM";
defparam ram_block1a30.operation_mode = "single_port";
defparam ram_block1a30.port_a_address_clear = "none";
defparam ram_block1a30.port_a_address_width = 13;
defparam ram_block1a30.port_a_byte_enable_mask_width = 1;
defparam ram_block1a30.port_a_byte_size = 1;
defparam ram_block1a30.port_a_data_out_clear = "none";
defparam ram_block1a30.port_a_data_out_clock = "none";
defparam ram_block1a30.port_a_data_width = 1;
defparam ram_block1a30.port_a_first_address = 0;
defparam ram_block1a30.port_a_first_bit_number = 30;
defparam ram_block1a30.port_a_last_address = 5119;
defparam ram_block1a30.port_a_logical_ram_depth = 5120;
defparam ram_block1a30.port_a_logical_ram_width = 32;
defparam ram_block1a30.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a30.ram_block_type = "auto";
defparam ram_block1a30.mem_init2 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a30.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a30.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a7(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a7_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a7.clk0_core_clock_enable = "ena0";
defparam ram_block1a7.clk0_input_clock_enable = "ena0";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.init_file = "processor_onchip_mem.hex";
defparam ram_block1a7.init_file_layout = "port_a";
defparam ram_block1a7.logical_ram_name = "processor_onchip_mem:onchip_mem|altsyncram:the_altsyncram|altsyncram_02n1:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.operation_mode = "single_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 13;
defparam ram_block1a7.port_a_byte_enable_mask_width = 1;
defparam ram_block1a7.port_a_byte_size = 1;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 5119;
defparam ram_block1a7.port_a_logical_ram_depth = 5120;
defparam ram_block1a7.port_a_logical_ram_width = 32;
defparam ram_block1a7.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a7.ram_block_type = "auto";
defparam ram_block1a7.mem_init2 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a7.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a7.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a23(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[23]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a23_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a23.clk0_core_clock_enable = "ena0";
defparam ram_block1a23.clk0_input_clock_enable = "ena0";
defparam ram_block1a23.data_interleave_offset_in_bits = 1;
defparam ram_block1a23.data_interleave_width_in_bits = 1;
defparam ram_block1a23.init_file = "processor_onchip_mem.hex";
defparam ram_block1a23.init_file_layout = "port_a";
defparam ram_block1a23.logical_ram_name = "processor_onchip_mem:onchip_mem|altsyncram:the_altsyncram|altsyncram_02n1:auto_generated|ALTSYNCRAM";
defparam ram_block1a23.operation_mode = "single_port";
defparam ram_block1a23.port_a_address_clear = "none";
defparam ram_block1a23.port_a_address_width = 13;
defparam ram_block1a23.port_a_byte_enable_mask_width = 1;
defparam ram_block1a23.port_a_byte_size = 1;
defparam ram_block1a23.port_a_data_out_clear = "none";
defparam ram_block1a23.port_a_data_out_clock = "none";
defparam ram_block1a23.port_a_data_width = 1;
defparam ram_block1a23.port_a_first_address = 0;
defparam ram_block1a23.port_a_first_bit_number = 23;
defparam ram_block1a23.port_a_last_address = 5119;
defparam ram_block1a23.port_a_logical_ram_depth = 5120;
defparam ram_block1a23.port_a_logical_ram_width = 32;
defparam ram_block1a23.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a23.ram_block_type = "auto";
defparam ram_block1a23.mem_init2 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a23.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a23.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a15(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a15_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a15.clk0_core_clock_enable = "ena0";
defparam ram_block1a15.clk0_input_clock_enable = "ena0";
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.init_file = "processor_onchip_mem.hex";
defparam ram_block1a15.init_file_layout = "port_a";
defparam ram_block1a15.logical_ram_name = "processor_onchip_mem:onchip_mem|altsyncram:the_altsyncram|altsyncram_02n1:auto_generated|ALTSYNCRAM";
defparam ram_block1a15.operation_mode = "single_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 13;
defparam ram_block1a15.port_a_byte_enable_mask_width = 1;
defparam ram_block1a15.port_a_byte_size = 1;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 5119;
defparam ram_block1a15.port_a_logical_ram_depth = 5120;
defparam ram_block1a15.port_a_logical_ram_width = 32;
defparam ram_block1a15.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a15.ram_block_type = "auto";
defparam ram_block1a15.mem_init2 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a15.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a15.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a31(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[31]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a31_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a31.clk0_core_clock_enable = "ena0";
defparam ram_block1a31.clk0_input_clock_enable = "ena0";
defparam ram_block1a31.data_interleave_offset_in_bits = 1;
defparam ram_block1a31.data_interleave_width_in_bits = 1;
defparam ram_block1a31.init_file = "processor_onchip_mem.hex";
defparam ram_block1a31.init_file_layout = "port_a";
defparam ram_block1a31.logical_ram_name = "processor_onchip_mem:onchip_mem|altsyncram:the_altsyncram|altsyncram_02n1:auto_generated|ALTSYNCRAM";
defparam ram_block1a31.operation_mode = "single_port";
defparam ram_block1a31.port_a_address_clear = "none";
defparam ram_block1a31.port_a_address_width = 13;
defparam ram_block1a31.port_a_byte_enable_mask_width = 1;
defparam ram_block1a31.port_a_byte_size = 1;
defparam ram_block1a31.port_a_data_out_clear = "none";
defparam ram_block1a31.port_a_data_out_clock = "none";
defparam ram_block1a31.port_a_data_width = 1;
defparam ram_block1a31.port_a_first_address = 0;
defparam ram_block1a31.port_a_first_bit_number = 31;
defparam ram_block1a31.port_a_last_address = 5119;
defparam ram_block1a31.port_a_logical_ram_depth = 5120;
defparam ram_block1a31.port_a_logical_ram_width = 32;
defparam ram_block1a31.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a31.ram_block_type = "auto";
defparam ram_block1a31.mem_init2 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a31.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a31.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a11(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a11_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a11.clk0_core_clock_enable = "ena0";
defparam ram_block1a11.clk0_input_clock_enable = "ena0";
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.init_file = "processor_onchip_mem.hex";
defparam ram_block1a11.init_file_layout = "port_a";
defparam ram_block1a11.logical_ram_name = "processor_onchip_mem:onchip_mem|altsyncram:the_altsyncram|altsyncram_02n1:auto_generated|ALTSYNCRAM";
defparam ram_block1a11.operation_mode = "single_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 13;
defparam ram_block1a11.port_a_byte_enable_mask_width = 1;
defparam ram_block1a11.port_a_byte_size = 1;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 5119;
defparam ram_block1a11.port_a_logical_ram_depth = 5120;
defparam ram_block1a11.port_a_logical_ram_width = 32;
defparam ram_block1a11.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a11.ram_block_type = "auto";
defparam ram_block1a11.mem_init2 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a11.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a11.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a27(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[27]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a27_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a27.clk0_core_clock_enable = "ena0";
defparam ram_block1a27.clk0_input_clock_enable = "ena0";
defparam ram_block1a27.data_interleave_offset_in_bits = 1;
defparam ram_block1a27.data_interleave_width_in_bits = 1;
defparam ram_block1a27.init_file = "processor_onchip_mem.hex";
defparam ram_block1a27.init_file_layout = "port_a";
defparam ram_block1a27.logical_ram_name = "processor_onchip_mem:onchip_mem|altsyncram:the_altsyncram|altsyncram_02n1:auto_generated|ALTSYNCRAM";
defparam ram_block1a27.operation_mode = "single_port";
defparam ram_block1a27.port_a_address_clear = "none";
defparam ram_block1a27.port_a_address_width = 13;
defparam ram_block1a27.port_a_byte_enable_mask_width = 1;
defparam ram_block1a27.port_a_byte_size = 1;
defparam ram_block1a27.port_a_data_out_clear = "none";
defparam ram_block1a27.port_a_data_out_clock = "none";
defparam ram_block1a27.port_a_data_width = 1;
defparam ram_block1a27.port_a_first_address = 0;
defparam ram_block1a27.port_a_first_bit_number = 27;
defparam ram_block1a27.port_a_last_address = 5119;
defparam ram_block1a27.port_a_logical_ram_depth = 5120;
defparam ram_block1a27.port_a_logical_ram_width = 32;
defparam ram_block1a27.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a27.ram_block_type = "auto";
defparam ram_block1a27.mem_init2 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a27.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a27.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a10(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a10_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a10.clk0_core_clock_enable = "ena0";
defparam ram_block1a10.clk0_input_clock_enable = "ena0";
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.init_file = "processor_onchip_mem.hex";
defparam ram_block1a10.init_file_layout = "port_a";
defparam ram_block1a10.logical_ram_name = "processor_onchip_mem:onchip_mem|altsyncram:the_altsyncram|altsyncram_02n1:auto_generated|ALTSYNCRAM";
defparam ram_block1a10.operation_mode = "single_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 13;
defparam ram_block1a10.port_a_byte_enable_mask_width = 1;
defparam ram_block1a10.port_a_byte_size = 1;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 5119;
defparam ram_block1a10.port_a_logical_ram_depth = 5120;
defparam ram_block1a10.port_a_logical_ram_width = 32;
defparam ram_block1a10.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a10.ram_block_type = "auto";
defparam ram_block1a10.mem_init2 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a10.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a10.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a26(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[26]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a26_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a26.clk0_core_clock_enable = "ena0";
defparam ram_block1a26.clk0_input_clock_enable = "ena0";
defparam ram_block1a26.data_interleave_offset_in_bits = 1;
defparam ram_block1a26.data_interleave_width_in_bits = 1;
defparam ram_block1a26.init_file = "processor_onchip_mem.hex";
defparam ram_block1a26.init_file_layout = "port_a";
defparam ram_block1a26.logical_ram_name = "processor_onchip_mem:onchip_mem|altsyncram:the_altsyncram|altsyncram_02n1:auto_generated|ALTSYNCRAM";
defparam ram_block1a26.operation_mode = "single_port";
defparam ram_block1a26.port_a_address_clear = "none";
defparam ram_block1a26.port_a_address_width = 13;
defparam ram_block1a26.port_a_byte_enable_mask_width = 1;
defparam ram_block1a26.port_a_byte_size = 1;
defparam ram_block1a26.port_a_data_out_clear = "none";
defparam ram_block1a26.port_a_data_out_clock = "none";
defparam ram_block1a26.port_a_data_width = 1;
defparam ram_block1a26.port_a_first_address = 0;
defparam ram_block1a26.port_a_first_bit_number = 26;
defparam ram_block1a26.port_a_last_address = 5119;
defparam ram_block1a26.port_a_logical_ram_depth = 5120;
defparam ram_block1a26.port_a_logical_ram_width = 32;
defparam ram_block1a26.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a26.ram_block_type = "auto";
defparam ram_block1a26.mem_init2 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a26.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a26.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a25(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[25]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a25_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a25.clk0_core_clock_enable = "ena0";
defparam ram_block1a25.clk0_input_clock_enable = "ena0";
defparam ram_block1a25.data_interleave_offset_in_bits = 1;
defparam ram_block1a25.data_interleave_width_in_bits = 1;
defparam ram_block1a25.init_file = "processor_onchip_mem.hex";
defparam ram_block1a25.init_file_layout = "port_a";
defparam ram_block1a25.logical_ram_name = "processor_onchip_mem:onchip_mem|altsyncram:the_altsyncram|altsyncram_02n1:auto_generated|ALTSYNCRAM";
defparam ram_block1a25.operation_mode = "single_port";
defparam ram_block1a25.port_a_address_clear = "none";
defparam ram_block1a25.port_a_address_width = 13;
defparam ram_block1a25.port_a_byte_enable_mask_width = 1;
defparam ram_block1a25.port_a_byte_size = 1;
defparam ram_block1a25.port_a_data_out_clear = "none";
defparam ram_block1a25.port_a_data_out_clock = "none";
defparam ram_block1a25.port_a_data_width = 1;
defparam ram_block1a25.port_a_first_address = 0;
defparam ram_block1a25.port_a_first_bit_number = 25;
defparam ram_block1a25.port_a_last_address = 5119;
defparam ram_block1a25.port_a_logical_ram_depth = 5120;
defparam ram_block1a25.port_a_logical_ram_width = 32;
defparam ram_block1a25.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a25.ram_block_type = "auto";
defparam ram_block1a25.mem_init2 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a25.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a25.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a9(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a9_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a9.clk0_core_clock_enable = "ena0";
defparam ram_block1a9.clk0_input_clock_enable = "ena0";
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.init_file = "processor_onchip_mem.hex";
defparam ram_block1a9.init_file_layout = "port_a";
defparam ram_block1a9.logical_ram_name = "processor_onchip_mem:onchip_mem|altsyncram:the_altsyncram|altsyncram_02n1:auto_generated|ALTSYNCRAM";
defparam ram_block1a9.operation_mode = "single_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 13;
defparam ram_block1a9.port_a_byte_enable_mask_width = 1;
defparam ram_block1a9.port_a_byte_size = 1;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 5119;
defparam ram_block1a9.port_a_logical_ram_depth = 5120;
defparam ram_block1a9.port_a_logical_ram_width = 32;
defparam ram_block1a9.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a9.ram_block_type = "auto";
defparam ram_block1a9.mem_init2 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a9.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a9.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a3(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a3_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a3.clk0_core_clock_enable = "ena0";
defparam ram_block1a3.clk0_input_clock_enable = "ena0";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.init_file = "processor_onchip_mem.hex";
defparam ram_block1a3.init_file_layout = "port_a";
defparam ram_block1a3.logical_ram_name = "processor_onchip_mem:onchip_mem|altsyncram:the_altsyncram|altsyncram_02n1:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.operation_mode = "single_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 13;
defparam ram_block1a3.port_a_byte_enable_mask_width = 1;
defparam ram_block1a3.port_a_byte_size = 1;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 5119;
defparam ram_block1a3.port_a_logical_ram_depth = 5120;
defparam ram_block1a3.port_a_logical_ram_width = 32;
defparam ram_block1a3.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a3.ram_block_type = "auto";
defparam ram_block1a3.mem_init2 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a3.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a3.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a19(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[19]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a19_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a19.clk0_core_clock_enable = "ena0";
defparam ram_block1a19.clk0_input_clock_enable = "ena0";
defparam ram_block1a19.data_interleave_offset_in_bits = 1;
defparam ram_block1a19.data_interleave_width_in_bits = 1;
defparam ram_block1a19.init_file = "processor_onchip_mem.hex";
defparam ram_block1a19.init_file_layout = "port_a";
defparam ram_block1a19.logical_ram_name = "processor_onchip_mem:onchip_mem|altsyncram:the_altsyncram|altsyncram_02n1:auto_generated|ALTSYNCRAM";
defparam ram_block1a19.operation_mode = "single_port";
defparam ram_block1a19.port_a_address_clear = "none";
defparam ram_block1a19.port_a_address_width = 13;
defparam ram_block1a19.port_a_byte_enable_mask_width = 1;
defparam ram_block1a19.port_a_byte_size = 1;
defparam ram_block1a19.port_a_data_out_clear = "none";
defparam ram_block1a19.port_a_data_out_clock = "none";
defparam ram_block1a19.port_a_data_width = 1;
defparam ram_block1a19.port_a_first_address = 0;
defparam ram_block1a19.port_a_first_bit_number = 19;
defparam ram_block1a19.port_a_last_address = 5119;
defparam ram_block1a19.port_a_logical_ram_depth = 5120;
defparam ram_block1a19.port_a_logical_ram_width = 32;
defparam ram_block1a19.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a19.ram_block_type = "auto";
defparam ram_block1a19.mem_init2 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a19.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a19.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a2(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a2_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a2.clk0_core_clock_enable = "ena0";
defparam ram_block1a2.clk0_input_clock_enable = "ena0";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.init_file = "processor_onchip_mem.hex";
defparam ram_block1a2.init_file_layout = "port_a";
defparam ram_block1a2.logical_ram_name = "processor_onchip_mem:onchip_mem|altsyncram:the_altsyncram|altsyncram_02n1:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.operation_mode = "single_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 13;
defparam ram_block1a2.port_a_byte_enable_mask_width = 1;
defparam ram_block1a2.port_a_byte_size = 1;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 5119;
defparam ram_block1a2.port_a_logical_ram_depth = 5120;
defparam ram_block1a2.port_a_logical_ram_width = 32;
defparam ram_block1a2.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a2.ram_block_type = "auto";
defparam ram_block1a2.mem_init2 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a2.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a2.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a18(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[18]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a18_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a18.clk0_core_clock_enable = "ena0";
defparam ram_block1a18.clk0_input_clock_enable = "ena0";
defparam ram_block1a18.data_interleave_offset_in_bits = 1;
defparam ram_block1a18.data_interleave_width_in_bits = 1;
defparam ram_block1a18.init_file = "processor_onchip_mem.hex";
defparam ram_block1a18.init_file_layout = "port_a";
defparam ram_block1a18.logical_ram_name = "processor_onchip_mem:onchip_mem|altsyncram:the_altsyncram|altsyncram_02n1:auto_generated|ALTSYNCRAM";
defparam ram_block1a18.operation_mode = "single_port";
defparam ram_block1a18.port_a_address_clear = "none";
defparam ram_block1a18.port_a_address_width = 13;
defparam ram_block1a18.port_a_byte_enable_mask_width = 1;
defparam ram_block1a18.port_a_byte_size = 1;
defparam ram_block1a18.port_a_data_out_clear = "none";
defparam ram_block1a18.port_a_data_out_clock = "none";
defparam ram_block1a18.port_a_data_width = 1;
defparam ram_block1a18.port_a_first_address = 0;
defparam ram_block1a18.port_a_first_bit_number = 18;
defparam ram_block1a18.port_a_last_address = 5119;
defparam ram_block1a18.port_a_logical_ram_depth = 5120;
defparam ram_block1a18.port_a_logical_ram_width = 32;
defparam ram_block1a18.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a18.ram_block_type = "auto";
defparam ram_block1a18.mem_init2 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a18.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a18.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a1(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a1_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a1.clk0_core_clock_enable = "ena0";
defparam ram_block1a1.clk0_input_clock_enable = "ena0";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.init_file = "processor_onchip_mem.hex";
defparam ram_block1a1.init_file_layout = "port_a";
defparam ram_block1a1.logical_ram_name = "processor_onchip_mem:onchip_mem|altsyncram:the_altsyncram|altsyncram_02n1:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.operation_mode = "single_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 13;
defparam ram_block1a1.port_a_byte_enable_mask_width = 1;
defparam ram_block1a1.port_a_byte_size = 1;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 5119;
defparam ram_block1a1.port_a_logical_ram_depth = 5120;
defparam ram_block1a1.port_a_logical_ram_width = 32;
defparam ram_block1a1.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a1.ram_block_type = "auto";
defparam ram_block1a1.mem_init2 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a1.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a1.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a17(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[17]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a17_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a17.clk0_core_clock_enable = "ena0";
defparam ram_block1a17.clk0_input_clock_enable = "ena0";
defparam ram_block1a17.data_interleave_offset_in_bits = 1;
defparam ram_block1a17.data_interleave_width_in_bits = 1;
defparam ram_block1a17.init_file = "processor_onchip_mem.hex";
defparam ram_block1a17.init_file_layout = "port_a";
defparam ram_block1a17.logical_ram_name = "processor_onchip_mem:onchip_mem|altsyncram:the_altsyncram|altsyncram_02n1:auto_generated|ALTSYNCRAM";
defparam ram_block1a17.operation_mode = "single_port";
defparam ram_block1a17.port_a_address_clear = "none";
defparam ram_block1a17.port_a_address_width = 13;
defparam ram_block1a17.port_a_byte_enable_mask_width = 1;
defparam ram_block1a17.port_a_byte_size = 1;
defparam ram_block1a17.port_a_data_out_clear = "none";
defparam ram_block1a17.port_a_data_out_clock = "none";
defparam ram_block1a17.port_a_data_width = 1;
defparam ram_block1a17.port_a_first_address = 0;
defparam ram_block1a17.port_a_first_bit_number = 17;
defparam ram_block1a17.port_a_last_address = 5119;
defparam ram_block1a17.port_a_logical_ram_depth = 5120;
defparam ram_block1a17.port_a_logical_ram_width = 32;
defparam ram_block1a17.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a17.ram_block_type = "auto";
defparam ram_block1a17.mem_init2 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a17.mem_init1 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
defparam ram_block1a17.mem_init0 = "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

endmodule

module processor_processor_switches_pio (
	r_sync_rst,
	M_alu_result_3,
	M_alu_result_2,
	readdata_0,
	readdata_8,
	readdata_5,
	readdata_4,
	readdata_6,
	readdata_7,
	readdata_9,
	readdata_3,
	readdata_2,
	readdata_1,
	clk_clk,
	switches_pio_external_connection_export_0,
	switches_pio_external_connection_export_8,
	switches_pio_external_connection_export_5,
	switches_pio_external_connection_export_4,
	switches_pio_external_connection_export_6,
	switches_pio_external_connection_export_7,
	switches_pio_external_connection_export_9,
	switches_pio_external_connection_export_3,
	switches_pio_external_connection_export_2,
	switches_pio_external_connection_export_1)/* synthesis synthesis_greybox=1 */;
input 	r_sync_rst;
input 	M_alu_result_3;
input 	M_alu_result_2;
output 	readdata_0;
output 	readdata_8;
output 	readdata_5;
output 	readdata_4;
output 	readdata_6;
output 	readdata_7;
output 	readdata_9;
output 	readdata_3;
output 	readdata_2;
output 	readdata_1;
input 	clk_clk;
input 	switches_pio_external_connection_export_0;
input 	switches_pio_external_connection_export_8;
input 	switches_pio_external_connection_export_5;
input 	switches_pio_external_connection_export_4;
input 	switches_pio_external_connection_export_6;
input 	switches_pio_external_connection_export_7;
input 	switches_pio_external_connection_export_9;
input 	switches_pio_external_connection_export_3;
input 	switches_pio_external_connection_export_2;
input 	switches_pio_external_connection_export_1;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \read_mux_out[0]~combout ;
wire \read_mux_out[8]~combout ;
wire \read_mux_out[5]~combout ;
wire \read_mux_out[4]~combout ;
wire \read_mux_out[6]~combout ;
wire \read_mux_out[7]~combout ;
wire \read_mux_out[9]~combout ;
wire \read_mux_out[3]~combout ;
wire \read_mux_out[2]~combout ;
wire \read_mux_out[1]~combout ;


dffeas \readdata[0] (
	.clk(clk_clk),
	.d(\read_mux_out[0]~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_0),
	.prn(vcc));
defparam \readdata[0] .is_wysiwyg = "true";
defparam \readdata[0] .power_up = "low";

dffeas \readdata[8] (
	.clk(clk_clk),
	.d(\read_mux_out[8]~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_8),
	.prn(vcc));
defparam \readdata[8] .is_wysiwyg = "true";
defparam \readdata[8] .power_up = "low";

dffeas \readdata[5] (
	.clk(clk_clk),
	.d(\read_mux_out[5]~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_5),
	.prn(vcc));
defparam \readdata[5] .is_wysiwyg = "true";
defparam \readdata[5] .power_up = "low";

dffeas \readdata[4] (
	.clk(clk_clk),
	.d(\read_mux_out[4]~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_4),
	.prn(vcc));
defparam \readdata[4] .is_wysiwyg = "true";
defparam \readdata[4] .power_up = "low";

dffeas \readdata[6] (
	.clk(clk_clk),
	.d(\read_mux_out[6]~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_6),
	.prn(vcc));
defparam \readdata[6] .is_wysiwyg = "true";
defparam \readdata[6] .power_up = "low";

dffeas \readdata[7] (
	.clk(clk_clk),
	.d(\read_mux_out[7]~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_7),
	.prn(vcc));
defparam \readdata[7] .is_wysiwyg = "true";
defparam \readdata[7] .power_up = "low";

dffeas \readdata[9] (
	.clk(clk_clk),
	.d(\read_mux_out[9]~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_9),
	.prn(vcc));
defparam \readdata[9] .is_wysiwyg = "true";
defparam \readdata[9] .power_up = "low";

dffeas \readdata[3] (
	.clk(clk_clk),
	.d(\read_mux_out[3]~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_3),
	.prn(vcc));
defparam \readdata[3] .is_wysiwyg = "true";
defparam \readdata[3] .power_up = "low";

dffeas \readdata[2] (
	.clk(clk_clk),
	.d(\read_mux_out[2]~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_2),
	.prn(vcc));
defparam \readdata[2] .is_wysiwyg = "true";
defparam \readdata[2] .power_up = "low";

dffeas \readdata[1] (
	.clk(clk_clk),
	.d(\read_mux_out[1]~combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_1),
	.prn(vcc));
defparam \readdata[1] .is_wysiwyg = "true";
defparam \readdata[1] .power_up = "low";

cyclonev_lcell_comb \read_mux_out[0] (
	.dataa(!M_alu_result_3),
	.datab(!M_alu_result_2),
	.datac(!switches_pio_external_connection_export_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[0]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[0] .extended_lut = "off";
defparam \read_mux_out[0] .lut_mask = 64'hEFEFEFEFEFEFEFEF;
defparam \read_mux_out[0] .shared_arith = "off";

cyclonev_lcell_comb \read_mux_out[8] (
	.dataa(!M_alu_result_3),
	.datab(!M_alu_result_2),
	.datac(!switches_pio_external_connection_export_8),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[8]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[8] .extended_lut = "off";
defparam \read_mux_out[8] .lut_mask = 64'hEFEFEFEFEFEFEFEF;
defparam \read_mux_out[8] .shared_arith = "off";

cyclonev_lcell_comb \read_mux_out[5] (
	.dataa(!M_alu_result_3),
	.datab(!M_alu_result_2),
	.datac(!switches_pio_external_connection_export_5),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[5]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[5] .extended_lut = "off";
defparam \read_mux_out[5] .lut_mask = 64'hEFEFEFEFEFEFEFEF;
defparam \read_mux_out[5] .shared_arith = "off";

cyclonev_lcell_comb \read_mux_out[4] (
	.dataa(!M_alu_result_3),
	.datab(!M_alu_result_2),
	.datac(!switches_pio_external_connection_export_4),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[4]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[4] .extended_lut = "off";
defparam \read_mux_out[4] .lut_mask = 64'hEFEFEFEFEFEFEFEF;
defparam \read_mux_out[4] .shared_arith = "off";

cyclonev_lcell_comb \read_mux_out[6] (
	.dataa(!M_alu_result_3),
	.datab(!M_alu_result_2),
	.datac(!switches_pio_external_connection_export_6),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[6]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[6] .extended_lut = "off";
defparam \read_mux_out[6] .lut_mask = 64'hEFEFEFEFEFEFEFEF;
defparam \read_mux_out[6] .shared_arith = "off";

cyclonev_lcell_comb \read_mux_out[7] (
	.dataa(!M_alu_result_3),
	.datab(!M_alu_result_2),
	.datac(!switches_pio_external_connection_export_7),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[7]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[7] .extended_lut = "off";
defparam \read_mux_out[7] .lut_mask = 64'hEFEFEFEFEFEFEFEF;
defparam \read_mux_out[7] .shared_arith = "off";

cyclonev_lcell_comb \read_mux_out[9] (
	.dataa(!M_alu_result_3),
	.datab(!M_alu_result_2),
	.datac(!switches_pio_external_connection_export_9),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[9]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[9] .extended_lut = "off";
defparam \read_mux_out[9] .lut_mask = 64'hEFEFEFEFEFEFEFEF;
defparam \read_mux_out[9] .shared_arith = "off";

cyclonev_lcell_comb \read_mux_out[3] (
	.dataa(!M_alu_result_3),
	.datab(!M_alu_result_2),
	.datac(!switches_pio_external_connection_export_3),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[3]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[3] .extended_lut = "off";
defparam \read_mux_out[3] .lut_mask = 64'hEFEFEFEFEFEFEFEF;
defparam \read_mux_out[3] .shared_arith = "off";

cyclonev_lcell_comb \read_mux_out[2] (
	.dataa(!M_alu_result_3),
	.datab(!M_alu_result_2),
	.datac(!switches_pio_external_connection_export_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[2]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[2] .extended_lut = "off";
defparam \read_mux_out[2] .lut_mask = 64'hEFEFEFEFEFEFEFEF;
defparam \read_mux_out[2] .shared_arith = "off";

cyclonev_lcell_comb \read_mux_out[1] (
	.dataa(!M_alu_result_3),
	.datab(!M_alu_result_2),
	.datac(!switches_pio_external_connection_export_1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[1]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[1] .extended_lut = "off";
defparam \read_mux_out[1] .lut_mask = 64'hEFEFEFEFEFEFEFEF;
defparam \read_mux_out[1] .shared_arith = "off";

endmodule

module processor_processor_sys_clk_timer (
	writedata,
	reset_n,
	clr_break_line,
	d_write,
	M_alu_result_5,
	M_alu_result_4,
	M_alu_result_6,
	Equal1,
	Equal2,
	M_alu_result_3,
	M_alu_result_2,
	mem_used_1,
	wait_latency_counter_1,
	wait_latency_counter_0,
	period_l_wr_strobe1,
	timeout_occurred1,
	control_register_0,
	readdata_0,
	readdata_8,
	readdata_5,
	readdata_13,
	readdata_4,
	readdata_12,
	readdata_6,
	readdata_14,
	readdata_7,
	readdata_15,
	readdata_11,
	readdata_10,
	readdata_9,
	readdata_3,
	readdata_2,
	readdata_1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	[15:0] writedata;
input 	reset_n;
input 	clr_break_line;
input 	d_write;
input 	M_alu_result_5;
input 	M_alu_result_4;
input 	M_alu_result_6;
input 	Equal1;
input 	Equal2;
input 	M_alu_result_3;
input 	M_alu_result_2;
input 	mem_used_1;
input 	wait_latency_counter_1;
input 	wait_latency_counter_0;
output 	period_l_wr_strobe1;
output 	timeout_occurred1;
output 	control_register_0;
output 	readdata_0;
output 	readdata_8;
output 	readdata_5;
output 	readdata_13;
output 	readdata_4;
output 	readdata_12;
output 	readdata_6;
output 	readdata_14;
output 	readdata_7;
output 	readdata_15;
output 	readdata_11;
output 	readdata_10;
output 	readdata_9;
output 	readdata_3;
output 	readdata_2;
output 	readdata_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \period_l_wr_strobe~1_combout ;
wire \status_wr_strobe~0_combout ;
wire \period_l_register[15]~4_combout ;
wire \Equal6~1_combout ;
wire \period_l_wr_strobe~combout ;
wire \period_l_register[15]~q ;
wire \period_l_register[3]~6_combout ;
wire \period_l_register[3]~q ;
wire \period_l_register[2]~7_combout ;
wire \period_l_register[2]~q ;
wire \period_l_register[1]~8_combout ;
wire \period_l_register[1]~q ;
wire \period_l_register[0]~0_combout ;
wire \period_l_register[0]~q ;
wire \Add0~113_sumout ;
wire \internal_counter~8_combout ;
wire \control_wr_strobe~combout ;
wire \control_register[1]~q ;
wire \force_reload~0_combout ;
wire \force_reload~q ;
wire \counter_is_running~0_combout ;
wire \counter_is_running~1_combout ;
wire \counter_is_running~q ;
wire \always0~1_combout ;
wire \internal_counter[0]~q ;
wire \Add0~114 ;
wire \Add0~109_sumout ;
wire \internal_counter~7_combout ;
wire \internal_counter[1]~q ;
wire \Add0~110 ;
wire \Add0~105_sumout ;
wire \internal_counter~6_combout ;
wire \internal_counter[2]~q ;
wire \Add0~106 ;
wire \Add0~101_sumout ;
wire \internal_counter~5_combout ;
wire \internal_counter[3]~q ;
wire \Add0~102 ;
wire \Add0~21_sumout ;
wire \period_l_register[4]~q ;
wire \internal_counter[4]~q ;
wire \period_l_register[9]~5_combout ;
wire \period_l_register[9]~q ;
wire \period_l_register[8]~1_combout ;
wire \period_l_register[8]~q ;
wire \period_l_register[6]~2_combout ;
wire \period_l_register[6]~q ;
wire \Add0~22 ;
wire \Add0~117_sumout ;
wire \period_l_register[5]~q ;
wire \internal_counter[5]~q ;
wire \Add0~118 ;
wire \Add0~97_sumout ;
wire \internal_counter~4_combout ;
wire \internal_counter[6]~q ;
wire \Add0~98 ;
wire \Add0~121_sumout ;
wire \period_l_register[7]~q ;
wire \internal_counter[7]~q ;
wire \Add0~122 ;
wire \Add0~93_sumout ;
wire \internal_counter~3_combout ;
wire \internal_counter[8]~q ;
wire \Add0~94 ;
wire \Add0~89_sumout ;
wire \internal_counter~2_combout ;
wire \internal_counter[9]~q ;
wire \Add0~90 ;
wire \Add0~125_sumout ;
wire \period_l_register[10]~q ;
wire \internal_counter[10]~q ;
wire \Add0~126 ;
wire \Add0~57_sumout ;
wire \period_l_register[11]~q ;
wire \internal_counter[11]~q ;
wire \Add0~58 ;
wire \Add0~61_sumout ;
wire \period_l_register[12]~q ;
wire \internal_counter[12]~q ;
wire \Add0~62 ;
wire \Add0~29_sumout ;
wire \period_l_register[13]~q ;
wire \internal_counter[13]~q ;
wire \Equal0~1_combout ;
wire \Equal0~2_combout ;
wire \Equal0~3_combout ;
wire \period_l_register[14]~3_combout ;
wire \period_l_register[14]~q ;
wire \Add0~30 ;
wire \Add0~85_sumout ;
wire \internal_counter~1_combout ;
wire \internal_counter[14]~q ;
wire \Equal0~4_combout ;
wire \Equal0~7_combout ;
wire \Equal0~8_combout ;
wire \always0~0_combout ;
wire \Add0~86 ;
wire \Add0~81_sumout ;
wire \internal_counter~0_combout ;
wire \internal_counter[15]~q ;
wire \Add0~82 ;
wire \Add0~25_sumout ;
wire \Equal6~0_combout ;
wire \period_h_wr_strobe~combout ;
wire \period_h_register[0]~q ;
wire \internal_counter[16]~q ;
wire \Add0~26 ;
wire \Add0~49_sumout ;
wire \period_h_register[1]~q ;
wire \internal_counter[17]~q ;
wire \Add0~50 ;
wire \Add0~77_sumout ;
wire \period_h_register[2]~q ;
wire \internal_counter[18]~q ;
wire \Add0~78 ;
wire \Add0~65_sumout ;
wire \period_h_register[3]~q ;
wire \internal_counter[19]~q ;
wire \Add0~66 ;
wire \Add0~33_sumout ;
wire \period_h_register[4]~q ;
wire \internal_counter[20]~q ;
wire \Add0~34 ;
wire \Add0~69_sumout ;
wire \period_h_register[5]~q ;
wire \internal_counter[21]~q ;
wire \Add0~70 ;
wire \Add0~73_sumout ;
wire \period_h_register[6]~q ;
wire \internal_counter[22]~q ;
wire \Add0~74 ;
wire \Add0~37_sumout ;
wire \period_h_register[7]~q ;
wire \internal_counter[23]~q ;
wire \Add0~38 ;
wire \Add0~41_sumout ;
wire \period_h_register[8]~q ;
wire \internal_counter[24]~q ;
wire \Add0~42 ;
wire \Add0~45_sumout ;
wire \period_h_register[9]~q ;
wire \internal_counter[25]~q ;
wire \Add0~46 ;
wire \Add0~5_sumout ;
wire \period_h_register[10]~q ;
wire \internal_counter[26]~q ;
wire \Add0~6 ;
wire \Add0~53_sumout ;
wire \period_h_register[11]~q ;
wire \internal_counter[27]~q ;
wire \Add0~54 ;
wire \Add0~9_sumout ;
wire \period_h_register[12]~q ;
wire \internal_counter[28]~q ;
wire \Add0~10 ;
wire \Add0~13_sumout ;
wire \period_h_register[13]~q ;
wire \internal_counter[29]~q ;
wire \Add0~14 ;
wire \Add0~17_sumout ;
wire \period_h_register[14]~q ;
wire \internal_counter[30]~q ;
wire \Add0~18 ;
wire \Add0~1_sumout ;
wire \period_h_register[15]~q ;
wire \internal_counter[31]~q ;
wire \Equal0~0_combout ;
wire \Equal0~5_combout ;
wire \Equal0~6_combout ;
wire \delayed_unxcounter_is_zeroxx0~q ;
wire \timeout_occurred~0_combout ;
wire \counter_snapshot[0]~0_combout ;
wire \snap_strobe~0_combout ;
wire \counter_snapshot[0]~q ;
wire \Equal6~2_combout ;
wire \read_mux_out[0]~0_combout ;
wire \counter_snapshot[16]~q ;
wire \read_mux_out[0]~1_combout ;
wire \read_mux_out[0]~combout ;
wire \counter_snapshot[8]~1_combout ;
wire \counter_snapshot[8]~q ;
wire \counter_snapshot[24]~q ;
wire \read_mux_out[8]~52_combout ;
wire \counter_snapshot[5]~q ;
wire \counter_snapshot[21]~q ;
wire \read_mux_out[5]~48_combout ;
wire \counter_snapshot[13]~q ;
wire \counter_snapshot[29]~q ;
wire \read_mux_out[13]~44_combout ;
wire \counter_snapshot[4]~q ;
wire \counter_snapshot[20]~q ;
wire \read_mux_out[4]~40_combout ;
wire \counter_snapshot[12]~q ;
wire \counter_snapshot[28]~q ;
wire \read_mux_out[12]~36_combout ;
wire \counter_snapshot[6]~2_combout ;
wire \counter_snapshot[6]~q ;
wire \counter_snapshot[22]~q ;
wire \read_mux_out[6]~32_combout ;
wire \counter_snapshot[14]~3_combout ;
wire \counter_snapshot[14]~q ;
wire \counter_snapshot[30]~q ;
wire \read_mux_out[14]~28_combout ;
wire \counter_snapshot[7]~q ;
wire \counter_snapshot[23]~q ;
wire \read_mux_out[7]~24_combout ;
wire \counter_snapshot[15]~4_combout ;
wire \counter_snapshot[15]~q ;
wire \counter_snapshot[31]~q ;
wire \read_mux_out[15]~20_combout ;
wire \counter_snapshot[11]~q ;
wire \counter_snapshot[27]~q ;
wire \read_mux_out[11]~16_combout ;
wire \counter_snapshot[10]~q ;
wire \counter_snapshot[26]~q ;
wire \read_mux_out[10]~12_combout ;
wire \counter_snapshot[9]~5_combout ;
wire \counter_snapshot[9]~q ;
wire \counter_snapshot[25]~q ;
wire \read_mux_out[9]~8_combout ;
wire \counter_snapshot[3]~6_combout ;
wire \counter_snapshot[3]~q ;
wire \read_mux_out[3]~2_combout ;
wire \counter_snapshot[19]~q ;
wire \control_register[3]~q ;
wire \read_mux_out[3]~3_combout ;
wire \read_mux_out[3]~combout ;
wire \counter_snapshot[2]~7_combout ;
wire \counter_snapshot[2]~q ;
wire \read_mux_out[2]~4_combout ;
wire \counter_snapshot[18]~q ;
wire \control_register[2]~q ;
wire \read_mux_out[2]~5_combout ;
wire \read_mux_out[2]~combout ;
wire \counter_snapshot[1]~8_combout ;
wire \counter_snapshot[1]~q ;
wire \read_mux_out[1]~6_combout ;
wire \counter_snapshot[17]~q ;
wire \read_mux_out[1]~7_combout ;
wire \read_mux_out[1]~combout ;


cyclonev_lcell_comb \period_l_wr_strobe~0 (
	.dataa(!clr_break_line),
	.datab(!M_alu_result_5),
	.datac(!M_alu_result_6),
	.datad(!Equal1),
	.datae(!Equal2),
	.dataf(!mem_used_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(period_l_wr_strobe1),
	.sumout(),
	.cout(),
	.shareout());
defparam \period_l_wr_strobe~0 .extended_lut = "off";
defparam \period_l_wr_strobe~0 .lut_mask = 64'hFFFFFFFFFDFFFFFF;
defparam \period_l_wr_strobe~0 .shared_arith = "off";

dffeas timeout_occurred(
	.clk(clk),
	.d(\timeout_occurred~0_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(timeout_occurred1),
	.prn(vcc));
defparam timeout_occurred.is_wysiwyg = "true";
defparam timeout_occurred.power_up = "low";

dffeas \control_register[0] (
	.clk(clk),
	.d(writedata[0]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\control_wr_strobe~combout ),
	.q(control_register_0),
	.prn(vcc));
defparam \control_register[0] .is_wysiwyg = "true";
defparam \control_register[0] .power_up = "low";

dffeas \readdata[0] (
	.clk(clk),
	.d(\read_mux_out[0]~combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_0),
	.prn(vcc));
defparam \readdata[0] .is_wysiwyg = "true";
defparam \readdata[0] .power_up = "low";

dffeas \readdata[8] (
	.clk(clk),
	.d(\read_mux_out[8]~52_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_8),
	.prn(vcc));
defparam \readdata[8] .is_wysiwyg = "true";
defparam \readdata[8] .power_up = "low";

dffeas \readdata[5] (
	.clk(clk),
	.d(\read_mux_out[5]~48_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_5),
	.prn(vcc));
defparam \readdata[5] .is_wysiwyg = "true";
defparam \readdata[5] .power_up = "low";

dffeas \readdata[13] (
	.clk(clk),
	.d(\read_mux_out[13]~44_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_13),
	.prn(vcc));
defparam \readdata[13] .is_wysiwyg = "true";
defparam \readdata[13] .power_up = "low";

dffeas \readdata[4] (
	.clk(clk),
	.d(\read_mux_out[4]~40_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_4),
	.prn(vcc));
defparam \readdata[4] .is_wysiwyg = "true";
defparam \readdata[4] .power_up = "low";

dffeas \readdata[12] (
	.clk(clk),
	.d(\read_mux_out[12]~36_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_12),
	.prn(vcc));
defparam \readdata[12] .is_wysiwyg = "true";
defparam \readdata[12] .power_up = "low";

dffeas \readdata[6] (
	.clk(clk),
	.d(\read_mux_out[6]~32_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_6),
	.prn(vcc));
defparam \readdata[6] .is_wysiwyg = "true";
defparam \readdata[6] .power_up = "low";

dffeas \readdata[14] (
	.clk(clk),
	.d(\read_mux_out[14]~28_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_14),
	.prn(vcc));
defparam \readdata[14] .is_wysiwyg = "true";
defparam \readdata[14] .power_up = "low";

dffeas \readdata[7] (
	.clk(clk),
	.d(\read_mux_out[7]~24_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_7),
	.prn(vcc));
defparam \readdata[7] .is_wysiwyg = "true";
defparam \readdata[7] .power_up = "low";

dffeas \readdata[15] (
	.clk(clk),
	.d(\read_mux_out[15]~20_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_15),
	.prn(vcc));
defparam \readdata[15] .is_wysiwyg = "true";
defparam \readdata[15] .power_up = "low";

dffeas \readdata[11] (
	.clk(clk),
	.d(\read_mux_out[11]~16_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_11),
	.prn(vcc));
defparam \readdata[11] .is_wysiwyg = "true";
defparam \readdata[11] .power_up = "low";

dffeas \readdata[10] (
	.clk(clk),
	.d(\read_mux_out[10]~12_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_10),
	.prn(vcc));
defparam \readdata[10] .is_wysiwyg = "true";
defparam \readdata[10] .power_up = "low";

dffeas \readdata[9] (
	.clk(clk),
	.d(\read_mux_out[9]~8_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_9),
	.prn(vcc));
defparam \readdata[9] .is_wysiwyg = "true";
defparam \readdata[9] .power_up = "low";

dffeas \readdata[3] (
	.clk(clk),
	.d(\read_mux_out[3]~combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_3),
	.prn(vcc));
defparam \readdata[3] .is_wysiwyg = "true";
defparam \readdata[3] .power_up = "low";

dffeas \readdata[2] (
	.clk(clk),
	.d(\read_mux_out[2]~combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_2),
	.prn(vcc));
defparam \readdata[2] .is_wysiwyg = "true";
defparam \readdata[2] .power_up = "low";

dffeas \readdata[1] (
	.clk(clk),
	.d(\read_mux_out[1]~combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_1),
	.prn(vcc));
defparam \readdata[1] .is_wysiwyg = "true";
defparam \readdata[1] .power_up = "low";

cyclonev_lcell_comb \period_l_wr_strobe~1 (
	.dataa(!d_write),
	.datab(!wait_latency_counter_1),
	.datac(!wait_latency_counter_0),
	.datad(!period_l_wr_strobe1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\period_l_wr_strobe~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \period_l_wr_strobe~1 .extended_lut = "off";
defparam \period_l_wr_strobe~1 .lut_mask = 64'hFDFFFDFFFDFFFDFF;
defparam \period_l_wr_strobe~1 .shared_arith = "off";

cyclonev_lcell_comb \status_wr_strobe~0 (
	.dataa(!M_alu_result_3),
	.datab(!M_alu_result_2),
	.datac(!M_alu_result_4),
	.datad(!\period_l_wr_strobe~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\status_wr_strobe~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \status_wr_strobe~0 .extended_lut = "off";
defparam \status_wr_strobe~0 .lut_mask = 64'hFEFFFEFFFEFFFEFF;
defparam \status_wr_strobe~0 .shared_arith = "off";

cyclonev_lcell_comb \period_l_register[15]~4 (
	.dataa(!writedata[15]),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\period_l_register[15]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \period_l_register[15]~4 .extended_lut = "off";
defparam \period_l_register[15]~4 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \period_l_register[15]~4 .shared_arith = "off";

cyclonev_lcell_comb \Equal6~1 (
	.dataa(!M_alu_result_3),
	.datab(!M_alu_result_2),
	.datac(!M_alu_result_4),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal6~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal6~1 .extended_lut = "off";
defparam \Equal6~1 .lut_mask = 64'hFDFDFDFDFDFDFDFD;
defparam \Equal6~1 .shared_arith = "off";

cyclonev_lcell_comb period_l_wr_strobe(
	.dataa(!\period_l_wr_strobe~1_combout ),
	.datab(!\Equal6~1_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\period_l_wr_strobe~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam period_l_wr_strobe.extended_lut = "off";
defparam period_l_wr_strobe.lut_mask = 64'h7777777777777777;
defparam period_l_wr_strobe.shared_arith = "off";

dffeas \period_l_register[15] (
	.clk(clk),
	.d(\period_l_register[15]~4_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\period_l_wr_strobe~combout ),
	.q(\period_l_register[15]~q ),
	.prn(vcc));
defparam \period_l_register[15] .is_wysiwyg = "true";
defparam \period_l_register[15] .power_up = "low";

cyclonev_lcell_comb \period_l_register[3]~6 (
	.dataa(!writedata[3]),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\period_l_register[3]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \period_l_register[3]~6 .extended_lut = "off";
defparam \period_l_register[3]~6 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \period_l_register[3]~6 .shared_arith = "off";

dffeas \period_l_register[3] (
	.clk(clk),
	.d(\period_l_register[3]~6_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\period_l_wr_strobe~combout ),
	.q(\period_l_register[3]~q ),
	.prn(vcc));
defparam \period_l_register[3] .is_wysiwyg = "true";
defparam \period_l_register[3] .power_up = "low";

cyclonev_lcell_comb \period_l_register[2]~7 (
	.dataa(!writedata[2]),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\period_l_register[2]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \period_l_register[2]~7 .extended_lut = "off";
defparam \period_l_register[2]~7 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \period_l_register[2]~7 .shared_arith = "off";

dffeas \period_l_register[2] (
	.clk(clk),
	.d(\period_l_register[2]~7_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\period_l_wr_strobe~combout ),
	.q(\period_l_register[2]~q ),
	.prn(vcc));
defparam \period_l_register[2] .is_wysiwyg = "true";
defparam \period_l_register[2] .power_up = "low";

cyclonev_lcell_comb \period_l_register[1]~8 (
	.dataa(!writedata[1]),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\period_l_register[1]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \period_l_register[1]~8 .extended_lut = "off";
defparam \period_l_register[1]~8 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \period_l_register[1]~8 .shared_arith = "off";

dffeas \period_l_register[1] (
	.clk(clk),
	.d(\period_l_register[1]~8_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\period_l_wr_strobe~combout ),
	.q(\period_l_register[1]~q ),
	.prn(vcc));
defparam \period_l_register[1] .is_wysiwyg = "true";
defparam \period_l_register[1] .power_up = "low";

cyclonev_lcell_comb \period_l_register[0]~0 (
	.dataa(!writedata[0]),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\period_l_register[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \period_l_register[0]~0 .extended_lut = "off";
defparam \period_l_register[0]~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \period_l_register[0]~0 .shared_arith = "off";

dffeas \period_l_register[0] (
	.clk(clk),
	.d(\period_l_register[0]~0_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\period_l_wr_strobe~combout ),
	.q(\period_l_register[0]~q ),
	.prn(vcc));
defparam \period_l_register[0] .is_wysiwyg = "true";
defparam \period_l_register[0] .power_up = "low";

cyclonev_lcell_comb \Add0~113 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\internal_counter[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~113_sumout ),
	.cout(\Add0~114 ),
	.shareout());
defparam \Add0~113 .extended_lut = "off";
defparam \Add0~113 .lut_mask = 64'h000000000000FF00;
defparam \Add0~113 .shared_arith = "off";

cyclonev_lcell_comb \internal_counter~8 (
	.dataa(!\period_l_register[0]~q ),
	.datab(!\always0~0_combout ),
	.datac(!\Add0~113_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\internal_counter~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \internal_counter~8 .extended_lut = "off";
defparam \internal_counter~8 .lut_mask = 64'hD1D1D1D1D1D1D1D1;
defparam \internal_counter~8 .shared_arith = "off";

cyclonev_lcell_comb control_wr_strobe(
	.dataa(!M_alu_result_3),
	.datab(!M_alu_result_2),
	.datac(!M_alu_result_4),
	.datad(!\period_l_wr_strobe~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\control_wr_strobe~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam control_wr_strobe.extended_lut = "off";
defparam control_wr_strobe.lut_mask = 64'hFBFFFBFFFBFFFBFF;
defparam control_wr_strobe.shared_arith = "off";

dffeas \control_register[1] (
	.clk(clk),
	.d(writedata[1]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\control_wr_strobe~combout ),
	.q(\control_register[1]~q ),
	.prn(vcc));
defparam \control_register[1] .is_wysiwyg = "true";
defparam \control_register[1] .power_up = "low";

cyclonev_lcell_comb \force_reload~0 (
	.dataa(!M_alu_result_3),
	.datab(!M_alu_result_4),
	.datac(!\period_l_wr_strobe~1_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\force_reload~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \force_reload~0 .extended_lut = "off";
defparam \force_reload~0 .lut_mask = 64'hDFDFDFDFDFDFDFDF;
defparam \force_reload~0 .shared_arith = "off";

dffeas force_reload(
	.clk(clk),
	.d(\force_reload~0_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\force_reload~q ),
	.prn(vcc));
defparam force_reload.is_wysiwyg = "true";
defparam force_reload.power_up = "low";

cyclonev_lcell_comb \counter_is_running~0 (
	.dataa(!\Equal0~6_combout ),
	.datab(!\control_register[1]~q ),
	.datac(!\counter_is_running~q ),
	.datad(!\force_reload~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\counter_is_running~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \counter_is_running~0 .extended_lut = "off";
defparam \counter_is_running~0 .lut_mask = 64'hFFBFFFBFFFBFFFBF;
defparam \counter_is_running~0 .shared_arith = "off";

cyclonev_lcell_comb \counter_is_running~1 (
	.dataa(!writedata[2]),
	.datab(!writedata[3]),
	.datac(!\control_wr_strobe~combout ),
	.datad(!\counter_is_running~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\counter_is_running~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \counter_is_running~1 .extended_lut = "off";
defparam \counter_is_running~1 .lut_mask = 64'hC5FFC5FFC5FFC5FF;
defparam \counter_is_running~1 .shared_arith = "off";

dffeas counter_is_running(
	.clk(clk),
	.d(\counter_is_running~1_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\counter_is_running~q ),
	.prn(vcc));
defparam counter_is_running.is_wysiwyg = "true";
defparam counter_is_running.power_up = "low";

cyclonev_lcell_comb \always0~1 (
	.dataa(!\counter_is_running~q ),
	.datab(!\force_reload~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always0~1 .extended_lut = "off";
defparam \always0~1 .lut_mask = 64'h7777777777777777;
defparam \always0~1 .shared_arith = "off";

dffeas \internal_counter[0] (
	.clk(clk),
	.d(\internal_counter~8_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(\internal_counter[0]~q ),
	.prn(vcc));
defparam \internal_counter[0] .is_wysiwyg = "true";
defparam \internal_counter[0] .power_up = "low";

cyclonev_lcell_comb \Add0~109 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\internal_counter[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~114 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~109_sumout ),
	.cout(\Add0~110 ),
	.shareout());
defparam \Add0~109 .extended_lut = "off";
defparam \Add0~109 .lut_mask = 64'h000000000000FF00;
defparam \Add0~109 .shared_arith = "off";

cyclonev_lcell_comb \internal_counter~7 (
	.dataa(!\period_l_register[1]~q ),
	.datab(!\always0~0_combout ),
	.datac(!\Add0~109_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\internal_counter~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \internal_counter~7 .extended_lut = "off";
defparam \internal_counter~7 .lut_mask = 64'hD1D1D1D1D1D1D1D1;
defparam \internal_counter~7 .shared_arith = "off";

dffeas \internal_counter[1] (
	.clk(clk),
	.d(\internal_counter~7_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(\internal_counter[1]~q ),
	.prn(vcc));
defparam \internal_counter[1] .is_wysiwyg = "true";
defparam \internal_counter[1] .power_up = "low";

cyclonev_lcell_comb \Add0~105 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\internal_counter[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~110 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~105_sumout ),
	.cout(\Add0~106 ),
	.shareout());
defparam \Add0~105 .extended_lut = "off";
defparam \Add0~105 .lut_mask = 64'h000000000000FF00;
defparam \Add0~105 .shared_arith = "off";

cyclonev_lcell_comb \internal_counter~6 (
	.dataa(!\period_l_register[2]~q ),
	.datab(!\always0~0_combout ),
	.datac(!\Add0~105_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\internal_counter~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \internal_counter~6 .extended_lut = "off";
defparam \internal_counter~6 .lut_mask = 64'hD1D1D1D1D1D1D1D1;
defparam \internal_counter~6 .shared_arith = "off";

dffeas \internal_counter[2] (
	.clk(clk),
	.d(\internal_counter~6_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(\internal_counter[2]~q ),
	.prn(vcc));
defparam \internal_counter[2] .is_wysiwyg = "true";
defparam \internal_counter[2] .power_up = "low";

cyclonev_lcell_comb \Add0~101 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\internal_counter[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~106 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~101_sumout ),
	.cout(\Add0~102 ),
	.shareout());
defparam \Add0~101 .extended_lut = "off";
defparam \Add0~101 .lut_mask = 64'h000000000000FF00;
defparam \Add0~101 .shared_arith = "off";

cyclonev_lcell_comb \internal_counter~5 (
	.dataa(!\period_l_register[3]~q ),
	.datab(!\always0~0_combout ),
	.datac(!\Add0~101_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\internal_counter~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \internal_counter~5 .extended_lut = "off";
defparam \internal_counter~5 .lut_mask = 64'hD1D1D1D1D1D1D1D1;
defparam \internal_counter~5 .shared_arith = "off";

dffeas \internal_counter[3] (
	.clk(clk),
	.d(\internal_counter~5_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(\internal_counter[3]~q ),
	.prn(vcc));
defparam \internal_counter[3] .is_wysiwyg = "true";
defparam \internal_counter[3] .power_up = "low";

cyclonev_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\internal_counter[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~102 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout());
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h00000000000000FF;
defparam \Add0~21 .shared_arith = "off";

dffeas \period_l_register[4] (
	.clk(clk),
	.d(writedata[4]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\period_l_wr_strobe~combout ),
	.q(\period_l_register[4]~q ),
	.prn(vcc));
defparam \period_l_register[4] .is_wysiwyg = "true";
defparam \period_l_register[4] .power_up = "low";

dffeas \internal_counter[4] (
	.clk(clk),
	.d(\Add0~21_sumout ),
	.asdata(\period_l_register[4]~q ),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always0~0_combout ),
	.ena(\always0~1_combout ),
	.q(\internal_counter[4]~q ),
	.prn(vcc));
defparam \internal_counter[4] .is_wysiwyg = "true";
defparam \internal_counter[4] .power_up = "low";

cyclonev_lcell_comb \period_l_register[9]~5 (
	.dataa(!writedata[9]),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\period_l_register[9]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \period_l_register[9]~5 .extended_lut = "off";
defparam \period_l_register[9]~5 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \period_l_register[9]~5 .shared_arith = "off";

dffeas \period_l_register[9] (
	.clk(clk),
	.d(\period_l_register[9]~5_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\period_l_wr_strobe~combout ),
	.q(\period_l_register[9]~q ),
	.prn(vcc));
defparam \period_l_register[9] .is_wysiwyg = "true";
defparam \period_l_register[9] .power_up = "low";

cyclonev_lcell_comb \period_l_register[8]~1 (
	.dataa(!writedata[8]),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\period_l_register[8]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \period_l_register[8]~1 .extended_lut = "off";
defparam \period_l_register[8]~1 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \period_l_register[8]~1 .shared_arith = "off";

dffeas \period_l_register[8] (
	.clk(clk),
	.d(\period_l_register[8]~1_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\period_l_wr_strobe~combout ),
	.q(\period_l_register[8]~q ),
	.prn(vcc));
defparam \period_l_register[8] .is_wysiwyg = "true";
defparam \period_l_register[8] .power_up = "low";

cyclonev_lcell_comb \period_l_register[6]~2 (
	.dataa(!writedata[6]),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\period_l_register[6]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \period_l_register[6]~2 .extended_lut = "off";
defparam \period_l_register[6]~2 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \period_l_register[6]~2 .shared_arith = "off";

dffeas \period_l_register[6] (
	.clk(clk),
	.d(\period_l_register[6]~2_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\period_l_wr_strobe~combout ),
	.q(\period_l_register[6]~q ),
	.prn(vcc));
defparam \period_l_register[6] .is_wysiwyg = "true";
defparam \period_l_register[6] .power_up = "low";

cyclonev_lcell_comb \Add0~117 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\internal_counter[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~117_sumout ),
	.cout(\Add0~118 ),
	.shareout());
defparam \Add0~117 .extended_lut = "off";
defparam \Add0~117 .lut_mask = 64'h00000000000000FF;
defparam \Add0~117 .shared_arith = "off";

dffeas \period_l_register[5] (
	.clk(clk),
	.d(writedata[5]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\period_l_wr_strobe~combout ),
	.q(\period_l_register[5]~q ),
	.prn(vcc));
defparam \period_l_register[5] .is_wysiwyg = "true";
defparam \period_l_register[5] .power_up = "low";

dffeas \internal_counter[5] (
	.clk(clk),
	.d(\Add0~117_sumout ),
	.asdata(\period_l_register[5]~q ),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always0~0_combout ),
	.ena(\always0~1_combout ),
	.q(\internal_counter[5]~q ),
	.prn(vcc));
defparam \internal_counter[5] .is_wysiwyg = "true";
defparam \internal_counter[5] .power_up = "low";

cyclonev_lcell_comb \Add0~97 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\internal_counter[6]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~118 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~97_sumout ),
	.cout(\Add0~98 ),
	.shareout());
defparam \Add0~97 .extended_lut = "off";
defparam \Add0~97 .lut_mask = 64'h000000000000FF00;
defparam \Add0~97 .shared_arith = "off";

cyclonev_lcell_comb \internal_counter~4 (
	.dataa(!\period_l_register[6]~q ),
	.datab(!\always0~0_combout ),
	.datac(!\Add0~97_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\internal_counter~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \internal_counter~4 .extended_lut = "off";
defparam \internal_counter~4 .lut_mask = 64'hD1D1D1D1D1D1D1D1;
defparam \internal_counter~4 .shared_arith = "off";

dffeas \internal_counter[6] (
	.clk(clk),
	.d(\internal_counter~4_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(\internal_counter[6]~q ),
	.prn(vcc));
defparam \internal_counter[6] .is_wysiwyg = "true";
defparam \internal_counter[6] .power_up = "low";

cyclonev_lcell_comb \Add0~121 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\internal_counter[7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~98 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~121_sumout ),
	.cout(\Add0~122 ),
	.shareout());
defparam \Add0~121 .extended_lut = "off";
defparam \Add0~121 .lut_mask = 64'h00000000000000FF;
defparam \Add0~121 .shared_arith = "off";

dffeas \period_l_register[7] (
	.clk(clk),
	.d(writedata[7]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\period_l_wr_strobe~combout ),
	.q(\period_l_register[7]~q ),
	.prn(vcc));
defparam \period_l_register[7] .is_wysiwyg = "true";
defparam \period_l_register[7] .power_up = "low";

dffeas \internal_counter[7] (
	.clk(clk),
	.d(\Add0~121_sumout ),
	.asdata(\period_l_register[7]~q ),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always0~0_combout ),
	.ena(\always0~1_combout ),
	.q(\internal_counter[7]~q ),
	.prn(vcc));
defparam \internal_counter[7] .is_wysiwyg = "true";
defparam \internal_counter[7] .power_up = "low";

cyclonev_lcell_comb \Add0~93 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\internal_counter[8]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~122 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~93_sumout ),
	.cout(\Add0~94 ),
	.shareout());
defparam \Add0~93 .extended_lut = "off";
defparam \Add0~93 .lut_mask = 64'h000000000000FF00;
defparam \Add0~93 .shared_arith = "off";

cyclonev_lcell_comb \internal_counter~3 (
	.dataa(!\period_l_register[8]~q ),
	.datab(!\always0~0_combout ),
	.datac(!\Add0~93_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\internal_counter~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \internal_counter~3 .extended_lut = "off";
defparam \internal_counter~3 .lut_mask = 64'hD1D1D1D1D1D1D1D1;
defparam \internal_counter~3 .shared_arith = "off";

dffeas \internal_counter[8] (
	.clk(clk),
	.d(\internal_counter~3_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(\internal_counter[8]~q ),
	.prn(vcc));
defparam \internal_counter[8] .is_wysiwyg = "true";
defparam \internal_counter[8] .power_up = "low";

cyclonev_lcell_comb \Add0~89 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\internal_counter[9]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~94 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~89_sumout ),
	.cout(\Add0~90 ),
	.shareout());
defparam \Add0~89 .extended_lut = "off";
defparam \Add0~89 .lut_mask = 64'h000000000000FF00;
defparam \Add0~89 .shared_arith = "off";

cyclonev_lcell_comb \internal_counter~2 (
	.dataa(!\period_l_register[9]~q ),
	.datab(!\always0~0_combout ),
	.datac(!\Add0~89_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\internal_counter~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \internal_counter~2 .extended_lut = "off";
defparam \internal_counter~2 .lut_mask = 64'hD1D1D1D1D1D1D1D1;
defparam \internal_counter~2 .shared_arith = "off";

dffeas \internal_counter[9] (
	.clk(clk),
	.d(\internal_counter~2_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(\internal_counter[9]~q ),
	.prn(vcc));
defparam \internal_counter[9] .is_wysiwyg = "true";
defparam \internal_counter[9] .power_up = "low";

cyclonev_lcell_comb \Add0~125 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\internal_counter[10]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~90 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~125_sumout ),
	.cout(\Add0~126 ),
	.shareout());
defparam \Add0~125 .extended_lut = "off";
defparam \Add0~125 .lut_mask = 64'h00000000000000FF;
defparam \Add0~125 .shared_arith = "off";

dffeas \period_l_register[10] (
	.clk(clk),
	.d(writedata[10]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\period_l_wr_strobe~combout ),
	.q(\period_l_register[10]~q ),
	.prn(vcc));
defparam \period_l_register[10] .is_wysiwyg = "true";
defparam \period_l_register[10] .power_up = "low";

dffeas \internal_counter[10] (
	.clk(clk),
	.d(\Add0~125_sumout ),
	.asdata(\period_l_register[10]~q ),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always0~0_combout ),
	.ena(\always0~1_combout ),
	.q(\internal_counter[10]~q ),
	.prn(vcc));
defparam \internal_counter[10] .is_wysiwyg = "true";
defparam \internal_counter[10] .power_up = "low";

cyclonev_lcell_comb \Add0~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\internal_counter[11]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~126 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~57_sumout ),
	.cout(\Add0~58 ),
	.shareout());
defparam \Add0~57 .extended_lut = "off";
defparam \Add0~57 .lut_mask = 64'h00000000000000FF;
defparam \Add0~57 .shared_arith = "off";

dffeas \period_l_register[11] (
	.clk(clk),
	.d(writedata[11]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\period_l_wr_strobe~combout ),
	.q(\period_l_register[11]~q ),
	.prn(vcc));
defparam \period_l_register[11] .is_wysiwyg = "true";
defparam \period_l_register[11] .power_up = "low";

dffeas \internal_counter[11] (
	.clk(clk),
	.d(\Add0~57_sumout ),
	.asdata(\period_l_register[11]~q ),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always0~0_combout ),
	.ena(\always0~1_combout ),
	.q(\internal_counter[11]~q ),
	.prn(vcc));
defparam \internal_counter[11] .is_wysiwyg = "true";
defparam \internal_counter[11] .power_up = "low";

cyclonev_lcell_comb \Add0~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\internal_counter[12]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~58 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~61_sumout ),
	.cout(\Add0~62 ),
	.shareout());
defparam \Add0~61 .extended_lut = "off";
defparam \Add0~61 .lut_mask = 64'h00000000000000FF;
defparam \Add0~61 .shared_arith = "off";

dffeas \period_l_register[12] (
	.clk(clk),
	.d(writedata[12]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\period_l_wr_strobe~combout ),
	.q(\period_l_register[12]~q ),
	.prn(vcc));
defparam \period_l_register[12] .is_wysiwyg = "true";
defparam \period_l_register[12] .power_up = "low";

dffeas \internal_counter[12] (
	.clk(clk),
	.d(\Add0~61_sumout ),
	.asdata(\period_l_register[12]~q ),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always0~0_combout ),
	.ena(\always0~1_combout ),
	.q(\internal_counter[12]~q ),
	.prn(vcc));
defparam \internal_counter[12] .is_wysiwyg = "true";
defparam \internal_counter[12] .power_up = "low";

cyclonev_lcell_comb \Add0~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\internal_counter[13]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~62 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~29_sumout ),
	.cout(\Add0~30 ),
	.shareout());
defparam \Add0~29 .extended_lut = "off";
defparam \Add0~29 .lut_mask = 64'h00000000000000FF;
defparam \Add0~29 .shared_arith = "off";

dffeas \period_l_register[13] (
	.clk(clk),
	.d(writedata[13]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\period_l_wr_strobe~combout ),
	.q(\period_l_register[13]~q ),
	.prn(vcc));
defparam \period_l_register[13] .is_wysiwyg = "true";
defparam \period_l_register[13] .power_up = "low";

dffeas \internal_counter[13] (
	.clk(clk),
	.d(\Add0~29_sumout ),
	.asdata(\period_l_register[13]~q ),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always0~0_combout ),
	.ena(\always0~1_combout ),
	.q(\internal_counter[13]~q ),
	.prn(vcc));
defparam \internal_counter[13] .is_wysiwyg = "true";
defparam \internal_counter[13] .power_up = "low";

cyclonev_lcell_comb \Equal0~1 (
	.dataa(!\internal_counter[28]~q ),
	.datab(!\internal_counter[29]~q ),
	.datac(!\internal_counter[30]~q ),
	.datad(!\internal_counter[4]~q ),
	.datae(!\internal_counter[16]~q ),
	.dataf(!\internal_counter[13]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~1 .extended_lut = "off";
defparam \Equal0~1 .lut_mask = 64'hFFFFFFFFFFFFFFFE;
defparam \Equal0~1 .shared_arith = "off";

cyclonev_lcell_comb \Equal0~2 (
	.dataa(!\internal_counter[20]~q ),
	.datab(!\internal_counter[23]~q ),
	.datac(!\internal_counter[24]~q ),
	.datad(!\internal_counter[25]~q ),
	.datae(!\internal_counter[17]~q ),
	.dataf(!\internal_counter[27]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~2 .extended_lut = "off";
defparam \Equal0~2 .lut_mask = 64'hFFFFFFFFFFFFFFFE;
defparam \Equal0~2 .shared_arith = "off";

cyclonev_lcell_comb \Equal0~3 (
	.dataa(!\internal_counter[11]~q ),
	.datab(!\internal_counter[12]~q ),
	.datac(!\internal_counter[19]~q ),
	.datad(!\internal_counter[21]~q ),
	.datae(!\internal_counter[22]~q ),
	.dataf(!\internal_counter[18]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~3 .extended_lut = "off";
defparam \Equal0~3 .lut_mask = 64'hFFFFFFFFFFFFFFFE;
defparam \Equal0~3 .shared_arith = "off";

cyclonev_lcell_comb \period_l_register[14]~3 (
	.dataa(!writedata[14]),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\period_l_register[14]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \period_l_register[14]~3 .extended_lut = "off";
defparam \period_l_register[14]~3 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \period_l_register[14]~3 .shared_arith = "off";

dffeas \period_l_register[14] (
	.clk(clk),
	.d(\period_l_register[14]~3_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\period_l_wr_strobe~combout ),
	.q(\period_l_register[14]~q ),
	.prn(vcc));
defparam \period_l_register[14] .is_wysiwyg = "true";
defparam \period_l_register[14] .power_up = "low";

cyclonev_lcell_comb \Add0~85 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\internal_counter[14]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~85_sumout ),
	.cout(\Add0~86 ),
	.shareout());
defparam \Add0~85 .extended_lut = "off";
defparam \Add0~85 .lut_mask = 64'h000000000000FF00;
defparam \Add0~85 .shared_arith = "off";

cyclonev_lcell_comb \internal_counter~1 (
	.dataa(!\period_l_register[14]~q ),
	.datab(!\always0~0_combout ),
	.datac(!\Add0~85_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\internal_counter~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \internal_counter~1 .extended_lut = "off";
defparam \internal_counter~1 .lut_mask = 64'hD1D1D1D1D1D1D1D1;
defparam \internal_counter~1 .shared_arith = "off";

dffeas \internal_counter[14] (
	.clk(clk),
	.d(\internal_counter~1_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(\internal_counter[14]~q ),
	.prn(vcc));
defparam \internal_counter[14] .is_wysiwyg = "true";
defparam \internal_counter[14] .power_up = "low";

cyclonev_lcell_comb \Equal0~4 (
	.dataa(!\internal_counter[15]~q ),
	.datab(!\internal_counter[14]~q ),
	.datac(!\internal_counter[9]~q ),
	.datad(!\internal_counter[8]~q ),
	.datae(!\internal_counter[6]~q ),
	.dataf(!\internal_counter[3]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~4 .extended_lut = "off";
defparam \Equal0~4 .lut_mask = 64'h7FFFFFFFFFFFFFFF;
defparam \Equal0~4 .shared_arith = "off";

cyclonev_lcell_comb \Equal0~7 (
	.dataa(!\internal_counter[2]~q ),
	.datab(!\internal_counter[1]~q ),
	.datac(!\internal_counter[0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~7 .extended_lut = "off";
defparam \Equal0~7 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \Equal0~7 .shared_arith = "off";

cyclonev_lcell_comb \Equal0~8 (
	.dataa(!\internal_counter[5]~q ),
	.datab(!\internal_counter[7]~q ),
	.datac(!\internal_counter[10]~q ),
	.datad(!\Equal0~4_combout ),
	.datae(!\Equal0~7_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~8 .extended_lut = "off";
defparam \Equal0~8 .lut_mask = 64'hFEFFFFFFFEFFFFFF;
defparam \Equal0~8 .shared_arith = "off";

cyclonev_lcell_comb \always0~0 (
	.dataa(!\Equal0~0_combout ),
	.datab(!\Equal0~1_combout ),
	.datac(!\Equal0~2_combout ),
	.datad(!\Equal0~3_combout ),
	.datae(!\Equal0~8_combout ),
	.dataf(!\force_reload~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always0~0 .extended_lut = "off";
defparam \always0~0 .lut_mask = 64'h7FFFFFFFFFFFFFFF;
defparam \always0~0 .shared_arith = "off";

cyclonev_lcell_comb \Add0~81 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\internal_counter[15]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~86 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~81_sumout ),
	.cout(\Add0~82 ),
	.shareout());
defparam \Add0~81 .extended_lut = "off";
defparam \Add0~81 .lut_mask = 64'h000000000000FF00;
defparam \Add0~81 .shared_arith = "off";

cyclonev_lcell_comb \internal_counter~0 (
	.dataa(!\period_l_register[15]~q ),
	.datab(!\always0~0_combout ),
	.datac(!\Add0~81_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\internal_counter~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \internal_counter~0 .extended_lut = "off";
defparam \internal_counter~0 .lut_mask = 64'hD1D1D1D1D1D1D1D1;
defparam \internal_counter~0 .shared_arith = "off";

dffeas \internal_counter[15] (
	.clk(clk),
	.d(\internal_counter~0_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(\internal_counter[15]~q ),
	.prn(vcc));
defparam \internal_counter[15] .is_wysiwyg = "true";
defparam \internal_counter[15] .power_up = "low";

cyclonev_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\internal_counter[16]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~82 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout());
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h00000000000000FF;
defparam \Add0~25 .shared_arith = "off";

cyclonev_lcell_comb \Equal6~0 (
	.dataa(!M_alu_result_3),
	.datab(!M_alu_result_2),
	.datac(!M_alu_result_4),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal6~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal6~0 .extended_lut = "off";
defparam \Equal6~0 .lut_mask = 64'hF7F7F7F7F7F7F7F7;
defparam \Equal6~0 .shared_arith = "off";

cyclonev_lcell_comb period_h_wr_strobe(
	.dataa(!\period_l_wr_strobe~1_combout ),
	.datab(!\Equal6~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\period_h_wr_strobe~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam period_h_wr_strobe.extended_lut = "off";
defparam period_h_wr_strobe.lut_mask = 64'h7777777777777777;
defparam period_h_wr_strobe.shared_arith = "off";

dffeas \period_h_register[0] (
	.clk(clk),
	.d(writedata[0]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\period_h_wr_strobe~combout ),
	.q(\period_h_register[0]~q ),
	.prn(vcc));
defparam \period_h_register[0] .is_wysiwyg = "true";
defparam \period_h_register[0] .power_up = "low";

dffeas \internal_counter[16] (
	.clk(clk),
	.d(\Add0~25_sumout ),
	.asdata(\period_h_register[0]~q ),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always0~0_combout ),
	.ena(\always0~1_combout ),
	.q(\internal_counter[16]~q ),
	.prn(vcc));
defparam \internal_counter[16] .is_wysiwyg = "true";
defparam \internal_counter[16] .power_up = "low";

cyclonev_lcell_comb \Add0~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\internal_counter[17]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~49_sumout ),
	.cout(\Add0~50 ),
	.shareout());
defparam \Add0~49 .extended_lut = "off";
defparam \Add0~49 .lut_mask = 64'h00000000000000FF;
defparam \Add0~49 .shared_arith = "off";

dffeas \period_h_register[1] (
	.clk(clk),
	.d(writedata[1]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\period_h_wr_strobe~combout ),
	.q(\period_h_register[1]~q ),
	.prn(vcc));
defparam \period_h_register[1] .is_wysiwyg = "true";
defparam \period_h_register[1] .power_up = "low";

dffeas \internal_counter[17] (
	.clk(clk),
	.d(\Add0~49_sumout ),
	.asdata(\period_h_register[1]~q ),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always0~0_combout ),
	.ena(\always0~1_combout ),
	.q(\internal_counter[17]~q ),
	.prn(vcc));
defparam \internal_counter[17] .is_wysiwyg = "true";
defparam \internal_counter[17] .power_up = "low";

cyclonev_lcell_comb \Add0~77 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\internal_counter[18]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~50 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~77_sumout ),
	.cout(\Add0~78 ),
	.shareout());
defparam \Add0~77 .extended_lut = "off";
defparam \Add0~77 .lut_mask = 64'h00000000000000FF;
defparam \Add0~77 .shared_arith = "off";

dffeas \period_h_register[2] (
	.clk(clk),
	.d(writedata[2]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\period_h_wr_strobe~combout ),
	.q(\period_h_register[2]~q ),
	.prn(vcc));
defparam \period_h_register[2] .is_wysiwyg = "true";
defparam \period_h_register[2] .power_up = "low";

dffeas \internal_counter[18] (
	.clk(clk),
	.d(\Add0~77_sumout ),
	.asdata(\period_h_register[2]~q ),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always0~0_combout ),
	.ena(\always0~1_combout ),
	.q(\internal_counter[18]~q ),
	.prn(vcc));
defparam \internal_counter[18] .is_wysiwyg = "true";
defparam \internal_counter[18] .power_up = "low";

cyclonev_lcell_comb \Add0~65 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\internal_counter[19]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~78 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~65_sumout ),
	.cout(\Add0~66 ),
	.shareout());
defparam \Add0~65 .extended_lut = "off";
defparam \Add0~65 .lut_mask = 64'h00000000000000FF;
defparam \Add0~65 .shared_arith = "off";

dffeas \period_h_register[3] (
	.clk(clk),
	.d(writedata[3]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\period_h_wr_strobe~combout ),
	.q(\period_h_register[3]~q ),
	.prn(vcc));
defparam \period_h_register[3] .is_wysiwyg = "true";
defparam \period_h_register[3] .power_up = "low";

dffeas \internal_counter[19] (
	.clk(clk),
	.d(\Add0~65_sumout ),
	.asdata(\period_h_register[3]~q ),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always0~0_combout ),
	.ena(\always0~1_combout ),
	.q(\internal_counter[19]~q ),
	.prn(vcc));
defparam \internal_counter[19] .is_wysiwyg = "true";
defparam \internal_counter[19] .power_up = "low";

cyclonev_lcell_comb \Add0~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\internal_counter[20]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~66 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~33_sumout ),
	.cout(\Add0~34 ),
	.shareout());
defparam \Add0~33 .extended_lut = "off";
defparam \Add0~33 .lut_mask = 64'h00000000000000FF;
defparam \Add0~33 .shared_arith = "off";

dffeas \period_h_register[4] (
	.clk(clk),
	.d(writedata[4]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\period_h_wr_strobe~combout ),
	.q(\period_h_register[4]~q ),
	.prn(vcc));
defparam \period_h_register[4] .is_wysiwyg = "true";
defparam \period_h_register[4] .power_up = "low";

dffeas \internal_counter[20] (
	.clk(clk),
	.d(\Add0~33_sumout ),
	.asdata(\period_h_register[4]~q ),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always0~0_combout ),
	.ena(\always0~1_combout ),
	.q(\internal_counter[20]~q ),
	.prn(vcc));
defparam \internal_counter[20] .is_wysiwyg = "true";
defparam \internal_counter[20] .power_up = "low";

cyclonev_lcell_comb \Add0~69 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\internal_counter[21]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~69_sumout ),
	.cout(\Add0~70 ),
	.shareout());
defparam \Add0~69 .extended_lut = "off";
defparam \Add0~69 .lut_mask = 64'h00000000000000FF;
defparam \Add0~69 .shared_arith = "off";

dffeas \period_h_register[5] (
	.clk(clk),
	.d(writedata[5]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\period_h_wr_strobe~combout ),
	.q(\period_h_register[5]~q ),
	.prn(vcc));
defparam \period_h_register[5] .is_wysiwyg = "true";
defparam \period_h_register[5] .power_up = "low";

dffeas \internal_counter[21] (
	.clk(clk),
	.d(\Add0~69_sumout ),
	.asdata(\period_h_register[5]~q ),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always0~0_combout ),
	.ena(\always0~1_combout ),
	.q(\internal_counter[21]~q ),
	.prn(vcc));
defparam \internal_counter[21] .is_wysiwyg = "true";
defparam \internal_counter[21] .power_up = "low";

cyclonev_lcell_comb \Add0~73 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\internal_counter[22]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~70 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~73_sumout ),
	.cout(\Add0~74 ),
	.shareout());
defparam \Add0~73 .extended_lut = "off";
defparam \Add0~73 .lut_mask = 64'h00000000000000FF;
defparam \Add0~73 .shared_arith = "off";

dffeas \period_h_register[6] (
	.clk(clk),
	.d(writedata[6]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\period_h_wr_strobe~combout ),
	.q(\period_h_register[6]~q ),
	.prn(vcc));
defparam \period_h_register[6] .is_wysiwyg = "true";
defparam \period_h_register[6] .power_up = "low";

dffeas \internal_counter[22] (
	.clk(clk),
	.d(\Add0~73_sumout ),
	.asdata(\period_h_register[6]~q ),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always0~0_combout ),
	.ena(\always0~1_combout ),
	.q(\internal_counter[22]~q ),
	.prn(vcc));
defparam \internal_counter[22] .is_wysiwyg = "true";
defparam \internal_counter[22] .power_up = "low";

cyclonev_lcell_comb \Add0~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\internal_counter[23]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~74 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~37_sumout ),
	.cout(\Add0~38 ),
	.shareout());
defparam \Add0~37 .extended_lut = "off";
defparam \Add0~37 .lut_mask = 64'h00000000000000FF;
defparam \Add0~37 .shared_arith = "off";

dffeas \period_h_register[7] (
	.clk(clk),
	.d(writedata[7]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\period_h_wr_strobe~combout ),
	.q(\period_h_register[7]~q ),
	.prn(vcc));
defparam \period_h_register[7] .is_wysiwyg = "true";
defparam \period_h_register[7] .power_up = "low";

dffeas \internal_counter[23] (
	.clk(clk),
	.d(\Add0~37_sumout ),
	.asdata(\period_h_register[7]~q ),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always0~0_combout ),
	.ena(\always0~1_combout ),
	.q(\internal_counter[23]~q ),
	.prn(vcc));
defparam \internal_counter[23] .is_wysiwyg = "true";
defparam \internal_counter[23] .power_up = "low";

cyclonev_lcell_comb \Add0~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\internal_counter[24]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~41_sumout ),
	.cout(\Add0~42 ),
	.shareout());
defparam \Add0~41 .extended_lut = "off";
defparam \Add0~41 .lut_mask = 64'h00000000000000FF;
defparam \Add0~41 .shared_arith = "off";

dffeas \period_h_register[8] (
	.clk(clk),
	.d(writedata[8]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\period_h_wr_strobe~combout ),
	.q(\period_h_register[8]~q ),
	.prn(vcc));
defparam \period_h_register[8] .is_wysiwyg = "true";
defparam \period_h_register[8] .power_up = "low";

dffeas \internal_counter[24] (
	.clk(clk),
	.d(\Add0~41_sumout ),
	.asdata(\period_h_register[8]~q ),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always0~0_combout ),
	.ena(\always0~1_combout ),
	.q(\internal_counter[24]~q ),
	.prn(vcc));
defparam \internal_counter[24] .is_wysiwyg = "true";
defparam \internal_counter[24] .power_up = "low";

cyclonev_lcell_comb \Add0~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\internal_counter[25]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~42 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~45_sumout ),
	.cout(\Add0~46 ),
	.shareout());
defparam \Add0~45 .extended_lut = "off";
defparam \Add0~45 .lut_mask = 64'h00000000000000FF;
defparam \Add0~45 .shared_arith = "off";

dffeas \period_h_register[9] (
	.clk(clk),
	.d(writedata[9]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\period_h_wr_strobe~combout ),
	.q(\period_h_register[9]~q ),
	.prn(vcc));
defparam \period_h_register[9] .is_wysiwyg = "true";
defparam \period_h_register[9] .power_up = "low";

dffeas \internal_counter[25] (
	.clk(clk),
	.d(\Add0~45_sumout ),
	.asdata(\period_h_register[9]~q ),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always0~0_combout ),
	.ena(\always0~1_combout ),
	.q(\internal_counter[25]~q ),
	.prn(vcc));
defparam \internal_counter[25] .is_wysiwyg = "true";
defparam \internal_counter[25] .power_up = "low";

cyclonev_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\internal_counter[26]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~46 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout());
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h00000000000000FF;
defparam \Add0~5 .shared_arith = "off";

dffeas \period_h_register[10] (
	.clk(clk),
	.d(writedata[10]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\period_h_wr_strobe~combout ),
	.q(\period_h_register[10]~q ),
	.prn(vcc));
defparam \period_h_register[10] .is_wysiwyg = "true";
defparam \period_h_register[10] .power_up = "low";

dffeas \internal_counter[26] (
	.clk(clk),
	.d(\Add0~5_sumout ),
	.asdata(\period_h_register[10]~q ),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always0~0_combout ),
	.ena(\always0~1_combout ),
	.q(\internal_counter[26]~q ),
	.prn(vcc));
defparam \internal_counter[26] .is_wysiwyg = "true";
defparam \internal_counter[26] .power_up = "low";

cyclonev_lcell_comb \Add0~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\internal_counter[27]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~53_sumout ),
	.cout(\Add0~54 ),
	.shareout());
defparam \Add0~53 .extended_lut = "off";
defparam \Add0~53 .lut_mask = 64'h00000000000000FF;
defparam \Add0~53 .shared_arith = "off";

dffeas \period_h_register[11] (
	.clk(clk),
	.d(writedata[11]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\period_h_wr_strobe~combout ),
	.q(\period_h_register[11]~q ),
	.prn(vcc));
defparam \period_h_register[11] .is_wysiwyg = "true";
defparam \period_h_register[11] .power_up = "low";

dffeas \internal_counter[27] (
	.clk(clk),
	.d(\Add0~53_sumout ),
	.asdata(\period_h_register[11]~q ),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always0~0_combout ),
	.ena(\always0~1_combout ),
	.q(\internal_counter[27]~q ),
	.prn(vcc));
defparam \internal_counter[27] .is_wysiwyg = "true";
defparam \internal_counter[27] .power_up = "low";

cyclonev_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\internal_counter[28]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~54 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout());
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h00000000000000FF;
defparam \Add0~9 .shared_arith = "off";

dffeas \period_h_register[12] (
	.clk(clk),
	.d(writedata[12]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\period_h_wr_strobe~combout ),
	.q(\period_h_register[12]~q ),
	.prn(vcc));
defparam \period_h_register[12] .is_wysiwyg = "true";
defparam \period_h_register[12] .power_up = "low";

dffeas \internal_counter[28] (
	.clk(clk),
	.d(\Add0~9_sumout ),
	.asdata(\period_h_register[12]~q ),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always0~0_combout ),
	.ena(\always0~1_combout ),
	.q(\internal_counter[28]~q ),
	.prn(vcc));
defparam \internal_counter[28] .is_wysiwyg = "true";
defparam \internal_counter[28] .power_up = "low";

cyclonev_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\internal_counter[29]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout());
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h00000000000000FF;
defparam \Add0~13 .shared_arith = "off";

dffeas \period_h_register[13] (
	.clk(clk),
	.d(writedata[13]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\period_h_wr_strobe~combout ),
	.q(\period_h_register[13]~q ),
	.prn(vcc));
defparam \period_h_register[13] .is_wysiwyg = "true";
defparam \period_h_register[13] .power_up = "low";

dffeas \internal_counter[29] (
	.clk(clk),
	.d(\Add0~13_sumout ),
	.asdata(\period_h_register[13]~q ),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always0~0_combout ),
	.ena(\always0~1_combout ),
	.q(\internal_counter[29]~q ),
	.prn(vcc));
defparam \internal_counter[29] .is_wysiwyg = "true";
defparam \internal_counter[29] .power_up = "low";

cyclonev_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\internal_counter[30]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout());
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h00000000000000FF;
defparam \Add0~17 .shared_arith = "off";

dffeas \period_h_register[14] (
	.clk(clk),
	.d(writedata[14]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\period_h_wr_strobe~combout ),
	.q(\period_h_register[14]~q ),
	.prn(vcc));
defparam \period_h_register[14] .is_wysiwyg = "true";
defparam \period_h_register[14] .power_up = "low";

dffeas \internal_counter[30] (
	.clk(clk),
	.d(\Add0~17_sumout ),
	.asdata(\period_h_register[14]~q ),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always0~0_combout ),
	.ena(\always0~1_combout ),
	.q(\internal_counter[30]~q ),
	.prn(vcc));
defparam \internal_counter[30] .is_wysiwyg = "true";
defparam \internal_counter[30] .power_up = "low";

cyclonev_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\internal_counter[31]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h00000000000000FF;
defparam \Add0~1 .shared_arith = "off";

dffeas \period_h_register[15] (
	.clk(clk),
	.d(writedata[15]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\period_h_wr_strobe~combout ),
	.q(\period_h_register[15]~q ),
	.prn(vcc));
defparam \period_h_register[15] .is_wysiwyg = "true";
defparam \period_h_register[15] .power_up = "low";

dffeas \internal_counter[31] (
	.clk(clk),
	.d(\Add0~1_sumout ),
	.asdata(\period_h_register[15]~q ),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\always0~0_combout ),
	.ena(\always0~1_combout ),
	.q(\internal_counter[31]~q ),
	.prn(vcc));
defparam \internal_counter[31] .is_wysiwyg = "true";
defparam \internal_counter[31] .power_up = "low";

cyclonev_lcell_comb \Equal0~0 (
	.dataa(!\internal_counter[31]~q ),
	.datab(!\internal_counter[26]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~0 .extended_lut = "off";
defparam \Equal0~0 .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \Equal0~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal0~5 (
	.dataa(!\internal_counter[2]~q ),
	.datab(!\internal_counter[1]~q ),
	.datac(!\internal_counter[0]~q ),
	.datad(!\internal_counter[5]~q ),
	.datae(!\internal_counter[7]~q ),
	.dataf(!\internal_counter[10]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~5 .extended_lut = "off";
defparam \Equal0~5 .lut_mask = 64'hFFFFFFFFFFFFFF7F;
defparam \Equal0~5 .shared_arith = "off";

cyclonev_lcell_comb \Equal0~6 (
	.dataa(!\Equal0~0_combout ),
	.datab(!\Equal0~1_combout ),
	.datac(!\Equal0~2_combout ),
	.datad(!\Equal0~3_combout ),
	.datae(!\Equal0~4_combout ),
	.dataf(!\Equal0~5_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~6 .extended_lut = "off";
defparam \Equal0~6 .lut_mask = 64'h7FFFFFFFFFFFFFFF;
defparam \Equal0~6 .shared_arith = "off";

dffeas delayed_unxcounter_is_zeroxx0(
	.clk(clk),
	.d(\Equal0~6_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\delayed_unxcounter_is_zeroxx0~q ),
	.prn(vcc));
defparam delayed_unxcounter_is_zeroxx0.is_wysiwyg = "true";
defparam delayed_unxcounter_is_zeroxx0.power_up = "low";

cyclonev_lcell_comb \timeout_occurred~0 (
	.dataa(!timeout_occurred1),
	.datab(!\status_wr_strobe~0_combout ),
	.datac(!\delayed_unxcounter_is_zeroxx0~q ),
	.datad(!\Equal0~6_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\timeout_occurred~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \timeout_occurred~0 .extended_lut = "off";
defparam \timeout_occurred~0 .lut_mask = 64'hFDFFFDFFFDFFFDFF;
defparam \timeout_occurred~0 .shared_arith = "off";

cyclonev_lcell_comb \counter_snapshot[0]~0 (
	.dataa(!\internal_counter[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\counter_snapshot[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \counter_snapshot[0]~0 .extended_lut = "off";
defparam \counter_snapshot[0]~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \counter_snapshot[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \snap_strobe~0 (
	.dataa(!M_alu_result_3),
	.datab(!M_alu_result_4),
	.datac(!\period_l_wr_strobe~1_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\snap_strobe~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \snap_strobe~0 .extended_lut = "off";
defparam \snap_strobe~0 .lut_mask = 64'hBFBFBFBFBFBFBFBF;
defparam \snap_strobe~0 .shared_arith = "off";

dffeas \counter_snapshot[0] (
	.clk(clk),
	.d(\counter_snapshot[0]~0_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\snap_strobe~0_combout ),
	.q(\counter_snapshot[0]~q ),
	.prn(vcc));
defparam \counter_snapshot[0] .is_wysiwyg = "true";
defparam \counter_snapshot[0] .power_up = "low";

cyclonev_lcell_comb \Equal6~2 (
	.dataa(!M_alu_result_3),
	.datab(!M_alu_result_2),
	.datac(!M_alu_result_4),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal6~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal6~2 .extended_lut = "off";
defparam \Equal6~2 .lut_mask = 64'hEFEFEFEFEFEFEFEF;
defparam \Equal6~2 .shared_arith = "off";

cyclonev_lcell_comb \read_mux_out[0]~0 (
	.dataa(!\period_l_register[0]~q ),
	.datab(!\Equal6~1_combout ),
	.datac(!\counter_snapshot[0]~q ),
	.datad(!\Equal6~2_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[0]~0 .extended_lut = "off";
defparam \read_mux_out[0]~0 .lut_mask = 64'hBFFFBFFFBFFFBFFF;
defparam \read_mux_out[0]~0 .shared_arith = "off";

dffeas \counter_snapshot[16] (
	.clk(clk),
	.d(\internal_counter[16]~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\snap_strobe~0_combout ),
	.q(\counter_snapshot[16]~q ),
	.prn(vcc));
defparam \counter_snapshot[16] .is_wysiwyg = "true";
defparam \counter_snapshot[16] .power_up = "low";

cyclonev_lcell_comb \read_mux_out[0]~1 (
	.dataa(!M_alu_result_3),
	.datab(!M_alu_result_2),
	.datac(!M_alu_result_4),
	.datad(!timeout_occurred1),
	.datae(!control_register_0),
	.dataf(!\counter_snapshot[16]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[0]~1 .extended_lut = "off";
defparam \read_mux_out[0]~1 .lut_mask = 64'hBEFFFFFFFFFFFFFF;
defparam \read_mux_out[0]~1 .shared_arith = "off";

cyclonev_lcell_comb \read_mux_out[0] (
	.dataa(!\period_h_register[0]~q ),
	.datab(!\Equal6~0_combout ),
	.datac(!\read_mux_out[0]~0_combout ),
	.datad(!\read_mux_out[0]~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[0]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[0] .extended_lut = "off";
defparam \read_mux_out[0] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \read_mux_out[0] .shared_arith = "off";

cyclonev_lcell_comb \counter_snapshot[8]~1 (
	.dataa(!\internal_counter[8]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\counter_snapshot[8]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \counter_snapshot[8]~1 .extended_lut = "off";
defparam \counter_snapshot[8]~1 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \counter_snapshot[8]~1 .shared_arith = "off";

dffeas \counter_snapshot[8] (
	.clk(clk),
	.d(\counter_snapshot[8]~1_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\snap_strobe~0_combout ),
	.q(\counter_snapshot[8]~q ),
	.prn(vcc));
defparam \counter_snapshot[8] .is_wysiwyg = "true";
defparam \counter_snapshot[8] .power_up = "low";

dffeas \counter_snapshot[24] (
	.clk(clk),
	.d(\internal_counter[24]~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\snap_strobe~0_combout ),
	.q(\counter_snapshot[24]~q ),
	.prn(vcc));
defparam \counter_snapshot[24] .is_wysiwyg = "true";
defparam \counter_snapshot[24] .power_up = "low";

cyclonev_lcell_comb \read_mux_out[8]~52 (
	.dataa(!M_alu_result_2),
	.datab(!M_alu_result_3),
	.datac(!\counter_snapshot[8]~q ),
	.datad(!\counter_snapshot[24]~q ),
	.datae(!M_alu_result_4),
	.dataf(!\period_h_register[8]~q ),
	.datag(!\period_l_register[8]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[8]~52_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[8]~52 .extended_lut = "on";
defparam \read_mux_out[8]~52 .lut_mask = 64'hFF6FFFF6FF6FFFF6;
defparam \read_mux_out[8]~52 .shared_arith = "off";

dffeas \counter_snapshot[5] (
	.clk(clk),
	.d(\internal_counter[5]~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\snap_strobe~0_combout ),
	.q(\counter_snapshot[5]~q ),
	.prn(vcc));
defparam \counter_snapshot[5] .is_wysiwyg = "true";
defparam \counter_snapshot[5] .power_up = "low";

dffeas \counter_snapshot[21] (
	.clk(clk),
	.d(\internal_counter[21]~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\snap_strobe~0_combout ),
	.q(\counter_snapshot[21]~q ),
	.prn(vcc));
defparam \counter_snapshot[21] .is_wysiwyg = "true";
defparam \counter_snapshot[21] .power_up = "low";

cyclonev_lcell_comb \read_mux_out[5]~48 (
	.dataa(!M_alu_result_2),
	.datab(!M_alu_result_3),
	.datac(!\counter_snapshot[5]~q ),
	.datad(!\counter_snapshot[21]~q ),
	.datae(!M_alu_result_4),
	.dataf(!\period_h_register[5]~q ),
	.datag(!\period_l_register[5]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[5]~48_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[5]~48 .extended_lut = "on";
defparam \read_mux_out[5]~48 .lut_mask = 64'hFFF6FFF6FFF6FFF6;
defparam \read_mux_out[5]~48 .shared_arith = "off";

dffeas \counter_snapshot[13] (
	.clk(clk),
	.d(\internal_counter[13]~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\snap_strobe~0_combout ),
	.q(\counter_snapshot[13]~q ),
	.prn(vcc));
defparam \counter_snapshot[13] .is_wysiwyg = "true";
defparam \counter_snapshot[13] .power_up = "low";

dffeas \counter_snapshot[29] (
	.clk(clk),
	.d(\internal_counter[29]~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\snap_strobe~0_combout ),
	.q(\counter_snapshot[29]~q ),
	.prn(vcc));
defparam \counter_snapshot[29] .is_wysiwyg = "true";
defparam \counter_snapshot[29] .power_up = "low";

cyclonev_lcell_comb \read_mux_out[13]~44 (
	.dataa(!M_alu_result_2),
	.datab(!M_alu_result_3),
	.datac(!\counter_snapshot[13]~q ),
	.datad(!\counter_snapshot[29]~q ),
	.datae(!M_alu_result_4),
	.dataf(!\period_h_register[13]~q ),
	.datag(!\period_l_register[13]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[13]~44_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[13]~44 .extended_lut = "on";
defparam \read_mux_out[13]~44 .lut_mask = 64'hFFF6FFF6FFF6FFF6;
defparam \read_mux_out[13]~44 .shared_arith = "off";

dffeas \counter_snapshot[4] (
	.clk(clk),
	.d(\internal_counter[4]~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\snap_strobe~0_combout ),
	.q(\counter_snapshot[4]~q ),
	.prn(vcc));
defparam \counter_snapshot[4] .is_wysiwyg = "true";
defparam \counter_snapshot[4] .power_up = "low";

dffeas \counter_snapshot[20] (
	.clk(clk),
	.d(\internal_counter[20]~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\snap_strobe~0_combout ),
	.q(\counter_snapshot[20]~q ),
	.prn(vcc));
defparam \counter_snapshot[20] .is_wysiwyg = "true";
defparam \counter_snapshot[20] .power_up = "low";

cyclonev_lcell_comb \read_mux_out[4]~40 (
	.dataa(!M_alu_result_2),
	.datab(!M_alu_result_3),
	.datac(!\counter_snapshot[4]~q ),
	.datad(!\counter_snapshot[20]~q ),
	.datae(!M_alu_result_4),
	.dataf(!\period_h_register[4]~q ),
	.datag(!\period_l_register[4]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[4]~40_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[4]~40 .extended_lut = "on";
defparam \read_mux_out[4]~40 .lut_mask = 64'hFFF6FFF6FFF6FFF6;
defparam \read_mux_out[4]~40 .shared_arith = "off";

dffeas \counter_snapshot[12] (
	.clk(clk),
	.d(\internal_counter[12]~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\snap_strobe~0_combout ),
	.q(\counter_snapshot[12]~q ),
	.prn(vcc));
defparam \counter_snapshot[12] .is_wysiwyg = "true";
defparam \counter_snapshot[12] .power_up = "low";

dffeas \counter_snapshot[28] (
	.clk(clk),
	.d(\internal_counter[28]~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\snap_strobe~0_combout ),
	.q(\counter_snapshot[28]~q ),
	.prn(vcc));
defparam \counter_snapshot[28] .is_wysiwyg = "true";
defparam \counter_snapshot[28] .power_up = "low";

cyclonev_lcell_comb \read_mux_out[12]~36 (
	.dataa(!M_alu_result_2),
	.datab(!M_alu_result_3),
	.datac(!\counter_snapshot[12]~q ),
	.datad(!\counter_snapshot[28]~q ),
	.datae(!M_alu_result_4),
	.dataf(!\period_h_register[12]~q ),
	.datag(!\period_l_register[12]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[12]~36_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[12]~36 .extended_lut = "on";
defparam \read_mux_out[12]~36 .lut_mask = 64'hFFF6FFF6FFF6FFF6;
defparam \read_mux_out[12]~36 .shared_arith = "off";

cyclonev_lcell_comb \counter_snapshot[6]~2 (
	.dataa(!\internal_counter[6]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\counter_snapshot[6]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \counter_snapshot[6]~2 .extended_lut = "off";
defparam \counter_snapshot[6]~2 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \counter_snapshot[6]~2 .shared_arith = "off";

dffeas \counter_snapshot[6] (
	.clk(clk),
	.d(\counter_snapshot[6]~2_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\snap_strobe~0_combout ),
	.q(\counter_snapshot[6]~q ),
	.prn(vcc));
defparam \counter_snapshot[6] .is_wysiwyg = "true";
defparam \counter_snapshot[6] .power_up = "low";

dffeas \counter_snapshot[22] (
	.clk(clk),
	.d(\internal_counter[22]~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\snap_strobe~0_combout ),
	.q(\counter_snapshot[22]~q ),
	.prn(vcc));
defparam \counter_snapshot[22] .is_wysiwyg = "true";
defparam \counter_snapshot[22] .power_up = "low";

cyclonev_lcell_comb \read_mux_out[6]~32 (
	.dataa(!M_alu_result_2),
	.datab(!M_alu_result_3),
	.datac(!\counter_snapshot[6]~q ),
	.datad(!\counter_snapshot[22]~q ),
	.datae(!M_alu_result_4),
	.dataf(!\period_h_register[6]~q ),
	.datag(!\period_l_register[6]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[6]~32_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[6]~32 .extended_lut = "on";
defparam \read_mux_out[6]~32 .lut_mask = 64'hFF6FFFF6FF6FFFF6;
defparam \read_mux_out[6]~32 .shared_arith = "off";

cyclonev_lcell_comb \counter_snapshot[14]~3 (
	.dataa(!\internal_counter[14]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\counter_snapshot[14]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \counter_snapshot[14]~3 .extended_lut = "off";
defparam \counter_snapshot[14]~3 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \counter_snapshot[14]~3 .shared_arith = "off";

dffeas \counter_snapshot[14] (
	.clk(clk),
	.d(\counter_snapshot[14]~3_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\snap_strobe~0_combout ),
	.q(\counter_snapshot[14]~q ),
	.prn(vcc));
defparam \counter_snapshot[14] .is_wysiwyg = "true";
defparam \counter_snapshot[14] .power_up = "low";

dffeas \counter_snapshot[30] (
	.clk(clk),
	.d(\internal_counter[30]~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\snap_strobe~0_combout ),
	.q(\counter_snapshot[30]~q ),
	.prn(vcc));
defparam \counter_snapshot[30] .is_wysiwyg = "true";
defparam \counter_snapshot[30] .power_up = "low";

cyclonev_lcell_comb \read_mux_out[14]~28 (
	.dataa(!M_alu_result_2),
	.datab(!M_alu_result_3),
	.datac(!\counter_snapshot[14]~q ),
	.datad(!\counter_snapshot[30]~q ),
	.datae(!M_alu_result_4),
	.dataf(!\period_h_register[14]~q ),
	.datag(!\period_l_register[14]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[14]~28_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[14]~28 .extended_lut = "on";
defparam \read_mux_out[14]~28 .lut_mask = 64'hFF6FFFF6FF6FFFF6;
defparam \read_mux_out[14]~28 .shared_arith = "off";

dffeas \counter_snapshot[7] (
	.clk(clk),
	.d(\internal_counter[7]~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\snap_strobe~0_combout ),
	.q(\counter_snapshot[7]~q ),
	.prn(vcc));
defparam \counter_snapshot[7] .is_wysiwyg = "true";
defparam \counter_snapshot[7] .power_up = "low";

dffeas \counter_snapshot[23] (
	.clk(clk),
	.d(\internal_counter[23]~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\snap_strobe~0_combout ),
	.q(\counter_snapshot[23]~q ),
	.prn(vcc));
defparam \counter_snapshot[23] .is_wysiwyg = "true";
defparam \counter_snapshot[23] .power_up = "low";

cyclonev_lcell_comb \read_mux_out[7]~24 (
	.dataa(!M_alu_result_2),
	.datab(!M_alu_result_3),
	.datac(!\counter_snapshot[7]~q ),
	.datad(!\counter_snapshot[23]~q ),
	.datae(!M_alu_result_4),
	.dataf(!\period_h_register[7]~q ),
	.datag(!\period_l_register[7]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[7]~24_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[7]~24 .extended_lut = "on";
defparam \read_mux_out[7]~24 .lut_mask = 64'hFFF6FFF6FFF6FFF6;
defparam \read_mux_out[7]~24 .shared_arith = "off";

cyclonev_lcell_comb \counter_snapshot[15]~4 (
	.dataa(!\internal_counter[15]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\counter_snapshot[15]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \counter_snapshot[15]~4 .extended_lut = "off";
defparam \counter_snapshot[15]~4 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \counter_snapshot[15]~4 .shared_arith = "off";

dffeas \counter_snapshot[15] (
	.clk(clk),
	.d(\counter_snapshot[15]~4_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\snap_strobe~0_combout ),
	.q(\counter_snapshot[15]~q ),
	.prn(vcc));
defparam \counter_snapshot[15] .is_wysiwyg = "true";
defparam \counter_snapshot[15] .power_up = "low";

dffeas \counter_snapshot[31] (
	.clk(clk),
	.d(\internal_counter[31]~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\snap_strobe~0_combout ),
	.q(\counter_snapshot[31]~q ),
	.prn(vcc));
defparam \counter_snapshot[31] .is_wysiwyg = "true";
defparam \counter_snapshot[31] .power_up = "low";

cyclonev_lcell_comb \read_mux_out[15]~20 (
	.dataa(!M_alu_result_2),
	.datab(!M_alu_result_3),
	.datac(!\counter_snapshot[15]~q ),
	.datad(!\counter_snapshot[31]~q ),
	.datae(!M_alu_result_4),
	.dataf(!\period_h_register[15]~q ),
	.datag(!\period_l_register[15]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[15]~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[15]~20 .extended_lut = "on";
defparam \read_mux_out[15]~20 .lut_mask = 64'hFF6FFFF6FF6FFFF6;
defparam \read_mux_out[15]~20 .shared_arith = "off";

dffeas \counter_snapshot[11] (
	.clk(clk),
	.d(\internal_counter[11]~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\snap_strobe~0_combout ),
	.q(\counter_snapshot[11]~q ),
	.prn(vcc));
defparam \counter_snapshot[11] .is_wysiwyg = "true";
defparam \counter_snapshot[11] .power_up = "low";

dffeas \counter_snapshot[27] (
	.clk(clk),
	.d(\internal_counter[27]~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\snap_strobe~0_combout ),
	.q(\counter_snapshot[27]~q ),
	.prn(vcc));
defparam \counter_snapshot[27] .is_wysiwyg = "true";
defparam \counter_snapshot[27] .power_up = "low";

cyclonev_lcell_comb \read_mux_out[11]~16 (
	.dataa(!M_alu_result_2),
	.datab(!M_alu_result_3),
	.datac(!\counter_snapshot[11]~q ),
	.datad(!\counter_snapshot[27]~q ),
	.datae(!M_alu_result_4),
	.dataf(!\period_h_register[11]~q ),
	.datag(!\period_l_register[11]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[11]~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[11]~16 .extended_lut = "on";
defparam \read_mux_out[11]~16 .lut_mask = 64'hFFF6FFF6FFF6FFF6;
defparam \read_mux_out[11]~16 .shared_arith = "off";

dffeas \counter_snapshot[10] (
	.clk(clk),
	.d(\internal_counter[10]~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\snap_strobe~0_combout ),
	.q(\counter_snapshot[10]~q ),
	.prn(vcc));
defparam \counter_snapshot[10] .is_wysiwyg = "true";
defparam \counter_snapshot[10] .power_up = "low";

dffeas \counter_snapshot[26] (
	.clk(clk),
	.d(\internal_counter[26]~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\snap_strobe~0_combout ),
	.q(\counter_snapshot[26]~q ),
	.prn(vcc));
defparam \counter_snapshot[26] .is_wysiwyg = "true";
defparam \counter_snapshot[26] .power_up = "low";

cyclonev_lcell_comb \read_mux_out[10]~12 (
	.dataa(!M_alu_result_2),
	.datab(!M_alu_result_3),
	.datac(!\counter_snapshot[10]~q ),
	.datad(!\counter_snapshot[26]~q ),
	.datae(!M_alu_result_4),
	.dataf(!\period_h_register[10]~q ),
	.datag(!\period_l_register[10]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[10]~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[10]~12 .extended_lut = "on";
defparam \read_mux_out[10]~12 .lut_mask = 64'hFFF6FFF6FFF6FFF6;
defparam \read_mux_out[10]~12 .shared_arith = "off";

cyclonev_lcell_comb \counter_snapshot[9]~5 (
	.dataa(!\internal_counter[9]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\counter_snapshot[9]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \counter_snapshot[9]~5 .extended_lut = "off";
defparam \counter_snapshot[9]~5 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \counter_snapshot[9]~5 .shared_arith = "off";

dffeas \counter_snapshot[9] (
	.clk(clk),
	.d(\counter_snapshot[9]~5_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\snap_strobe~0_combout ),
	.q(\counter_snapshot[9]~q ),
	.prn(vcc));
defparam \counter_snapshot[9] .is_wysiwyg = "true";
defparam \counter_snapshot[9] .power_up = "low";

dffeas \counter_snapshot[25] (
	.clk(clk),
	.d(\internal_counter[25]~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\snap_strobe~0_combout ),
	.q(\counter_snapshot[25]~q ),
	.prn(vcc));
defparam \counter_snapshot[25] .is_wysiwyg = "true";
defparam \counter_snapshot[25] .power_up = "low";

cyclonev_lcell_comb \read_mux_out[9]~8 (
	.dataa(!M_alu_result_2),
	.datab(!M_alu_result_3),
	.datac(!\counter_snapshot[9]~q ),
	.datad(!\counter_snapshot[25]~q ),
	.datae(!M_alu_result_4),
	.dataf(!\period_h_register[9]~q ),
	.datag(!\period_l_register[9]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[9]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[9]~8 .extended_lut = "on";
defparam \read_mux_out[9]~8 .lut_mask = 64'hFF6FFFF6FF6FFFF6;
defparam \read_mux_out[9]~8 .shared_arith = "off";

cyclonev_lcell_comb \counter_snapshot[3]~6 (
	.dataa(!\internal_counter[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\counter_snapshot[3]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \counter_snapshot[3]~6 .extended_lut = "off";
defparam \counter_snapshot[3]~6 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \counter_snapshot[3]~6 .shared_arith = "off";

dffeas \counter_snapshot[3] (
	.clk(clk),
	.d(\counter_snapshot[3]~6_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\snap_strobe~0_combout ),
	.q(\counter_snapshot[3]~q ),
	.prn(vcc));
defparam \counter_snapshot[3] .is_wysiwyg = "true";
defparam \counter_snapshot[3] .power_up = "low";

cyclonev_lcell_comb \read_mux_out[3]~2 (
	.dataa(!\Equal6~1_combout ),
	.datab(!\Equal6~2_combout ),
	.datac(!\period_l_register[3]~q ),
	.datad(!\counter_snapshot[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[3]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[3]~2 .extended_lut = "off";
defparam \read_mux_out[3]~2 .lut_mask = 64'hF7FFF7FFF7FFF7FF;
defparam \read_mux_out[3]~2 .shared_arith = "off";

dffeas \counter_snapshot[19] (
	.clk(clk),
	.d(\internal_counter[19]~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\snap_strobe~0_combout ),
	.q(\counter_snapshot[19]~q ),
	.prn(vcc));
defparam \counter_snapshot[19] .is_wysiwyg = "true";
defparam \counter_snapshot[19] .power_up = "low";

dffeas \control_register[3] (
	.clk(clk),
	.d(writedata[3]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\control_wr_strobe~combout ),
	.q(\control_register[3]~q ),
	.prn(vcc));
defparam \control_register[3] .is_wysiwyg = "true";
defparam \control_register[3] .power_up = "low";

cyclonev_lcell_comb \read_mux_out[3]~3 (
	.dataa(!M_alu_result_3),
	.datab(!M_alu_result_2),
	.datac(!M_alu_result_4),
	.datad(!\counter_snapshot[19]~q ),
	.datae(!\control_register[3]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[3]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[3]~3 .extended_lut = "off";
defparam \read_mux_out[3]~3 .lut_mask = 64'hA3FFFFFFA3FFFFFF;
defparam \read_mux_out[3]~3 .shared_arith = "off";

cyclonev_lcell_comb \read_mux_out[3] (
	.dataa(!\Equal6~0_combout ),
	.datab(!\period_h_register[3]~q ),
	.datac(!\read_mux_out[3]~2_combout ),
	.datad(!\read_mux_out[3]~3_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[3]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[3] .extended_lut = "off";
defparam \read_mux_out[3] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \read_mux_out[3] .shared_arith = "off";

cyclonev_lcell_comb \counter_snapshot[2]~7 (
	.dataa(!\internal_counter[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\counter_snapshot[2]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \counter_snapshot[2]~7 .extended_lut = "off";
defparam \counter_snapshot[2]~7 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \counter_snapshot[2]~7 .shared_arith = "off";

dffeas \counter_snapshot[2] (
	.clk(clk),
	.d(\counter_snapshot[2]~7_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\snap_strobe~0_combout ),
	.q(\counter_snapshot[2]~q ),
	.prn(vcc));
defparam \counter_snapshot[2] .is_wysiwyg = "true";
defparam \counter_snapshot[2] .power_up = "low";

cyclonev_lcell_comb \read_mux_out[2]~4 (
	.dataa(!\Equal6~1_combout ),
	.datab(!\Equal6~2_combout ),
	.datac(!\period_l_register[2]~q ),
	.datad(!\counter_snapshot[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[2]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[2]~4 .extended_lut = "off";
defparam \read_mux_out[2]~4 .lut_mask = 64'hF7FFF7FFF7FFF7FF;
defparam \read_mux_out[2]~4 .shared_arith = "off";

dffeas \counter_snapshot[18] (
	.clk(clk),
	.d(\internal_counter[18]~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\snap_strobe~0_combout ),
	.q(\counter_snapshot[18]~q ),
	.prn(vcc));
defparam \counter_snapshot[18] .is_wysiwyg = "true";
defparam \counter_snapshot[18] .power_up = "low";

dffeas \control_register[2] (
	.clk(clk),
	.d(writedata[2]),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\control_wr_strobe~combout ),
	.q(\control_register[2]~q ),
	.prn(vcc));
defparam \control_register[2] .is_wysiwyg = "true";
defparam \control_register[2] .power_up = "low";

cyclonev_lcell_comb \read_mux_out[2]~5 (
	.dataa(!M_alu_result_3),
	.datab(!M_alu_result_2),
	.datac(!M_alu_result_4),
	.datad(!\counter_snapshot[18]~q ),
	.datae(!\control_register[2]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[2]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[2]~5 .extended_lut = "off";
defparam \read_mux_out[2]~5 .lut_mask = 64'hA3FFFFFFA3FFFFFF;
defparam \read_mux_out[2]~5 .shared_arith = "off";

cyclonev_lcell_comb \read_mux_out[2] (
	.dataa(!\Equal6~0_combout ),
	.datab(!\period_h_register[2]~q ),
	.datac(!\read_mux_out[2]~4_combout ),
	.datad(!\read_mux_out[2]~5_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[2]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[2] .extended_lut = "off";
defparam \read_mux_out[2] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \read_mux_out[2] .shared_arith = "off";

cyclonev_lcell_comb \counter_snapshot[1]~8 (
	.dataa(!\internal_counter[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\counter_snapshot[1]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \counter_snapshot[1]~8 .extended_lut = "off";
defparam \counter_snapshot[1]~8 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \counter_snapshot[1]~8 .shared_arith = "off";

dffeas \counter_snapshot[1] (
	.clk(clk),
	.d(\counter_snapshot[1]~8_combout ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\snap_strobe~0_combout ),
	.q(\counter_snapshot[1]~q ),
	.prn(vcc));
defparam \counter_snapshot[1] .is_wysiwyg = "true";
defparam \counter_snapshot[1] .power_up = "low";

cyclonev_lcell_comb \read_mux_out[1]~6 (
	.dataa(!\Equal6~1_combout ),
	.datab(!\Equal6~2_combout ),
	.datac(!\period_l_register[1]~q ),
	.datad(!\counter_snapshot[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[1]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[1]~6 .extended_lut = "off";
defparam \read_mux_out[1]~6 .lut_mask = 64'hF7FFF7FFF7FFF7FF;
defparam \read_mux_out[1]~6 .shared_arith = "off";

dffeas \counter_snapshot[17] (
	.clk(clk),
	.d(\internal_counter[17]~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\snap_strobe~0_combout ),
	.q(\counter_snapshot[17]~q ),
	.prn(vcc));
defparam \counter_snapshot[17] .is_wysiwyg = "true";
defparam \counter_snapshot[17] .power_up = "low";

cyclonev_lcell_comb \read_mux_out[1]~7 (
	.dataa(!M_alu_result_3),
	.datab(!M_alu_result_2),
	.datac(!M_alu_result_4),
	.datad(!\counter_snapshot[17]~q ),
	.datae(!\control_register[1]~q ),
	.dataf(!\counter_is_running~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[1]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[1]~7 .extended_lut = "off";
defparam \read_mux_out[1]~7 .lut_mask = 64'hBEFFFFFFFFFFFFFF;
defparam \read_mux_out[1]~7 .shared_arith = "off";

cyclonev_lcell_comb \read_mux_out[1] (
	.dataa(!\Equal6~0_combout ),
	.datab(!\period_h_register[1]~q ),
	.datac(!\read_mux_out[1]~6_combout ),
	.datad(!\read_mux_out[1]~7_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_mux_out[1]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_mux_out[1] .extended_lut = "off";
defparam \read_mux_out[1] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \read_mux_out[1] .shared_arith = "off";

endmodule
