module clockControl;
endmodule
